entity hello is
end;

architecture behav of hello is
begin
  assert false report "Hello";
end behav;
