package p is
  -- as functions are longer in definitions, it might be written before
  function log2(param : positive) return natural;
end p;


