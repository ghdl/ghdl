package bb is new work.b generic map ( X => 6);

