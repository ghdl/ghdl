use work.b.all;

package c is
    subtype a1 is bit;
    subtype a2 is bit;
    subtype a3 is bit;
    subtype a4 is bit;
    subtype a5 is bit;
    subtype a6 is bit;
    subtype a7 is bit;
    subtype a8 is bit;
    subtype a9 is bit;
    subtype a10 is bit;
    subtype a11 is bit;
    subtype a12 is bit;
    subtype a13 is bit;
    subtype a14 is bit;
    subtype a15 is bit;
    subtype a16 is bit;
    subtype a17 is bit;
    subtype a18 is bit;
    subtype a19 is bit;
    subtype a20 is bit;
    subtype a21 is bit;
    subtype a22 is bit;
    subtype a23 is bit;
    subtype a24 is bit;
    subtype a25 is bit;
    subtype a26 is bit;
    subtype a27 is bit;
    subtype a28 is bit;
    subtype a29 is bit;
    subtype a30 is bit;
    subtype a31 is bit;
    subtype a32 is bit;
    subtype a33 is bit;
    subtype a34 is bit;
    subtype a35 is bit;
    subtype a36 is bit;
    subtype a37 is bit;
    subtype a38 is bit;
    subtype a39 is bit;
    subtype a40 is bit;
    subtype a41 is bit;
    subtype a42 is bit;
    subtype a43 is bit;
    subtype a44 is bit;
    subtype a45 is bit;
    subtype a46 is bit;
    subtype a47 is bit;
    subtype a48 is bit;
    subtype a49 is bit;
    subtype a50 is bit;
    subtype a51 is bit;
    subtype a52 is bit;
    subtype a53 is bit;
    subtype a54 is bit;
    subtype a55 is bit;
    subtype a56 is bit;
    subtype a57 is bit;
    subtype a58 is bit;
    subtype a59 is bit;
    subtype a60 is bit;
    subtype a61 is bit;
    subtype a62 is bit;
    subtype a63 is bit;
    subtype a64 is bit;
    subtype a65 is bit;
    subtype a66 is bit;
    subtype a67 is bit;
    subtype a68 is bit;
    subtype a69 is bit;
    subtype a70 is bit;
    subtype a71 is bit;
    subtype a72 is bit;
    subtype a73 is bit;
    subtype a74 is bit;
    subtype a75 is bit;
    subtype a76 is bit;
    subtype a77 is bit;
    subtype a78 is bit;
    subtype a79 is bit;
    subtype a80 is bit;
    subtype a81 is bit;
    subtype a82 is bit;
    subtype a83 is bit;
    subtype a84 is bit;
    subtype a85 is bit;
    subtype a86 is bit;
    subtype a87 is bit;
    subtype a88 is bit;
    subtype a89 is bit;
    subtype a90 is bit;
    subtype a91 is bit;
    subtype a92 is bit;
    subtype a93 is bit;
    subtype a94 is bit;
    subtype a95 is bit;
    subtype a96 is bit;
    subtype a97 is bit;
    subtype a98 is bit;
    subtype a99 is bit;
    subtype a100 is bit;
    subtype a101 is bit;
    subtype a102 is bit;
    subtype a103 is bit;
    subtype a104 is bit;
    subtype a105 is bit;
    subtype a106 is bit;
    subtype a107 is bit;
    subtype a108 is bit;
    subtype a109 is bit;
    subtype a110 is bit;
    subtype a111 is bit;
    subtype a112 is bit;
    subtype a113 is bit;
    subtype a114 is bit;
    subtype a115 is bit;
    subtype a116 is bit;
    subtype a117 is bit;
    subtype a118 is bit;
    subtype a119 is bit;
    subtype a120 is bit;
    subtype a121 is bit;
    subtype a122 is bit;
    subtype a123 is bit;
    subtype a124 is bit;
    subtype a125 is bit;
    subtype a126 is bit;
    subtype a127 is bit;
    subtype a128 is bit;
    subtype a129 is bit;
    subtype a130 is bit;
    subtype a131 is bit;
    subtype a132 is bit;
    subtype a133 is bit;
    subtype a134 is bit;
    subtype a135 is bit;
    subtype a136 is bit;
    subtype a137 is bit;
    subtype a138 is bit;
    subtype a139 is bit;
    subtype a140 is bit;
    subtype a141 is bit;
    subtype a142 is bit;
    subtype a143 is bit;
    subtype a144 is bit;
    subtype a145 is bit;
    subtype a146 is bit;
    subtype a147 is bit;
    subtype a148 is bit;
    subtype a149 is bit;
    subtype a150 is bit;
    subtype a151 is bit;
    subtype a152 is bit;
    subtype a153 is bit;
    subtype a154 is bit;
    subtype a155 is bit;
    subtype a156 is bit;
    subtype a157 is bit;
    subtype a158 is bit;
    subtype a159 is bit;
    subtype a160 is bit;
    subtype a161 is bit;
    subtype a162 is bit;
    subtype a163 is bit;
    subtype a164 is bit;
    subtype a165 is bit;
    subtype a166 is bit;
    subtype a167 is bit;
    subtype a168 is bit;
    subtype a169 is bit;
    subtype a170 is bit;
    subtype a171 is bit;
    subtype a172 is bit;
    subtype a173 is bit;
    subtype a174 is bit;
    subtype a175 is bit;
    subtype a176 is bit;
    subtype a177 is bit;
    subtype a178 is bit;
    subtype a179 is bit;
    subtype a180 is bit;
    subtype a181 is bit;
    subtype a182 is bit;
    subtype a183 is bit;
    subtype a184 is bit;
    subtype a185 is bit;
    subtype a186 is bit;
    subtype a187 is bit;
    subtype a188 is bit;
    subtype a189 is bit;
    subtype a190 is bit;
    subtype a191 is bit;
    subtype a192 is bit;
    subtype a193 is bit;
    subtype a194 is bit;
    subtype a195 is bit;
    subtype a196 is bit;
    subtype a197 is bit;
    subtype a198 is bit;
    subtype a199 is bit;
    subtype a200 is bit;
    subtype a201 is bit;
    subtype a202 is bit;
    subtype a203 is bit;
    subtype a204 is bit;
    subtype a205 is bit;
    subtype a206 is bit;
    subtype a207 is bit;
    subtype a208 is bit;
    subtype a209 is bit;
    subtype a210 is bit;
    subtype a211 is bit;
    subtype a212 is bit;
    subtype a213 is bit;
    subtype a214 is bit;
    subtype a215 is bit;
    subtype a216 is bit;
    subtype a217 is bit;
    subtype a218 is bit;
    subtype a219 is bit;
    subtype a220 is bit;
    subtype a221 is bit;
    subtype a222 is bit;
    subtype a223 is bit;
    subtype a224 is bit;
    subtype a225 is bit;
    subtype a226 is bit;
    subtype a227 is bit;
    subtype a228 is bit;
    subtype a229 is bit;
    subtype a230 is bit;
    subtype a231 is bit;
    subtype a232 is bit;
    subtype a233 is bit;
    subtype a234 is bit;
    subtype a235 is bit;
    subtype a236 is bit;
    subtype a237 is bit;
    subtype a238 is bit;
    subtype a239 is bit;
    subtype a240 is bit;
    subtype a241 is bit;
    subtype a242 is bit;
    subtype a243 is bit;
    subtype a244 is bit;
    subtype a245 is bit;
    subtype a246 is bit;
    subtype a247 is bit;
    subtype a248 is bit;
    subtype a249 is bit;
    subtype a250 is bit;
    subtype a251 is bit;
    subtype a252 is bit;
    subtype a253 is bit;
    subtype a254 is bit;
    subtype a255 is bit;
    subtype a256 is bit;
    subtype a257 is bit;
    subtype a258 is bit;
    subtype a259 is bit;
    subtype a260 is bit;
    subtype a261 is bit;
    subtype a262 is bit;
    subtype a263 is bit;
    subtype a264 is bit;
    subtype a265 is bit;
    subtype a266 is bit;
    subtype a267 is bit;
    subtype a268 is bit;
    subtype a269 is bit;
    subtype a270 is bit;
    subtype a271 is bit;
    subtype a272 is bit;
    subtype a273 is bit;
    subtype a274 is bit;
    subtype a275 is bit;
    subtype a276 is bit;
    subtype a277 is bit;
    subtype a278 is bit;
    subtype a279 is bit;
    subtype a280 is bit;
    subtype a281 is bit;
    subtype a282 is bit;
    subtype a283 is bit;
    subtype a284 is bit;
    subtype a285 is bit;
    subtype a286 is bit;
    subtype a287 is bit;
    subtype a288 is bit;
    subtype a289 is bit;
    subtype a290 is bit;
    subtype a291 is bit;
    subtype a292 is bit;
    subtype a293 is bit;
    subtype a294 is bit;
    subtype a295 is bit;
    subtype a296 is bit;
    subtype a297 is bit;
    subtype a298 is bit;
    subtype a299 is bit;
    subtype a300 is bit;
    subtype a301 is bit;
    subtype a302 is bit;
    subtype a303 is bit;
    subtype a304 is bit;
    subtype a305 is bit;
    subtype a306 is bit;
    subtype a307 is bit;
    subtype a308 is bit;
    subtype a309 is bit;
    subtype a310 is bit;
    subtype a311 is bit;
    subtype a312 is bit;
    subtype a313 is bit;
    subtype a314 is bit;
    subtype a315 is bit;
    subtype a316 is bit;
    subtype a317 is bit;
    subtype a318 is bit;
    subtype a319 is bit;
    subtype a320 is bit;
    subtype a321 is bit;
    subtype a322 is bit;
    subtype a323 is bit;
    subtype a324 is bit;
    subtype a325 is bit;
    subtype a326 is bit;
    subtype a327 is bit;
    subtype a328 is bit;
    subtype a329 is bit;
    subtype a330 is bit;
    subtype a331 is bit;
    subtype a332 is bit;
    subtype a333 is bit;
    subtype a334 is bit;
    subtype a335 is bit;
    subtype a336 is bit;
    subtype a337 is bit;
    subtype a338 is bit;
    subtype a339 is bit;
    subtype a340 is bit;
    subtype a341 is bit;
    subtype a342 is bit;
    subtype a343 is bit;
    subtype a344 is bit;
    subtype a345 is bit;
    subtype a346 is bit;
    subtype a347 is bit;
    subtype a348 is bit;
    subtype a349 is bit;
    subtype a350 is bit;
    subtype a351 is bit;
    subtype a352 is bit;
    subtype a353 is bit;
    subtype a354 is bit;
    subtype a355 is bit;
    subtype a356 is bit;
    subtype a357 is bit;
    subtype a358 is bit;
    subtype a359 is bit;
    subtype a360 is bit;
    subtype a361 is bit;
    subtype a362 is bit;
    subtype a363 is bit;
    subtype a364 is bit;
    subtype a365 is bit;
    subtype a366 is bit;
    subtype a367 is bit;
    subtype a368 is bit;
    subtype a369 is bit;
    subtype a370 is bit;
    subtype a371 is bit;
    subtype a372 is bit;
    subtype a373 is bit;
    subtype a374 is bit;
    subtype a375 is bit;
    subtype a376 is bit;
    subtype a377 is bit;
    subtype a378 is bit;
    subtype a379 is bit;
    subtype a380 is bit;
    subtype a381 is bit;
    subtype a382 is bit;
    subtype a383 is bit;
    subtype a384 is bit;
    subtype a385 is bit;
    subtype a386 is bit;
    subtype a387 is bit;
    subtype a388 is bit;
    subtype a389 is bit;
    subtype a390 is bit;
    subtype a391 is bit;
    subtype a392 is bit;
    subtype a393 is bit;
    subtype a394 is bit;
    subtype a395 is bit;
    subtype a396 is bit;
    subtype a397 is bit;
    subtype a398 is bit;
    subtype a399 is bit;
    subtype a400 is bit;
    subtype a401 is bit;
    subtype a402 is bit;
    subtype a403 is bit;
    subtype a404 is bit;
    subtype a405 is bit;
    subtype a406 is bit;
    subtype a407 is bit;
    subtype a408 is bit;
    subtype a409 is bit;
    subtype a410 is bit;
    subtype a411 is bit;
    subtype a412 is bit;
    subtype a413 is bit;
    subtype a414 is bit;
    subtype a415 is bit;
    subtype a416 is bit;
    subtype a417 is bit;
    subtype a418 is bit;
    subtype a419 is bit;
    subtype a420 is bit;
    subtype a421 is bit;
    subtype a422 is bit;
    subtype a423 is bit;
    subtype a424 is bit;
    subtype a425 is bit;
    subtype a426 is bit;
    subtype a427 is bit;
    subtype a428 is bit;
    subtype a429 is bit;
    subtype a430 is bit;
    subtype a431 is bit;
    subtype a432 is bit;
    subtype a433 is bit;
    subtype a434 is bit;
    subtype a435 is bit;
    subtype a436 is bit;
    subtype a437 is bit;
    subtype a438 is bit;
    subtype a439 is bit;
    subtype a440 is bit;
    subtype a441 is bit;
    subtype a442 is bit;
    subtype a443 is bit;
    subtype a444 is bit;
    subtype a445 is bit;
    subtype a446 is bit;
    subtype a447 is bit;
    subtype a448 is bit;
    subtype a449 is bit;
    subtype a450 is bit;
    subtype a451 is bit;
    subtype a452 is bit;
    subtype a453 is bit;
    subtype a454 is bit;
    subtype a455 is bit;
    subtype a456 is bit;
    subtype a457 is bit;
    subtype a458 is bit;
    subtype a459 is bit;
    subtype a460 is bit;
    subtype a461 is bit;
    subtype a462 is bit;
    subtype a463 is bit;
    subtype a464 is bit;
    subtype a465 is bit;
    subtype a466 is bit;
    subtype a467 is bit;
    subtype a468 is bit;
    subtype a469 is bit;
    subtype a470 is bit;
    subtype a471 is bit;
    subtype a472 is bit;
    subtype a473 is bit;
    subtype a474 is bit;
    subtype a475 is bit;
    subtype a476 is bit;
    subtype a477 is bit;
    subtype a478 is bit;
    subtype a479 is bit;
    subtype a480 is bit;
    subtype a481 is bit;
    subtype a482 is bit;
    subtype a483 is bit;
    subtype a484 is bit;
    subtype a485 is bit;
    subtype a486 is bit;
    subtype a487 is bit;
    subtype a488 is bit;
    subtype a489 is bit;
    subtype a490 is bit;
    subtype a491 is bit;
    subtype a492 is bit;
    subtype a493 is bit;
    subtype a494 is bit;
    subtype a495 is bit;
    subtype a496 is bit;
    subtype a497 is bit;
    subtype a498 is bit;
    subtype a499 is bit;
    subtype a500 is bit;
    subtype a501 is bit;
    subtype a502 is bit;
    subtype a503 is bit;
    subtype a504 is bit;
    subtype a505 is bit;
    subtype a506 is bit;
    subtype a507 is bit;
    subtype a508 is bit;
    subtype a509 is bit;
    subtype a510 is bit;
    subtype a511 is bit;
    subtype a512 is bit;
    subtype a513 is bit;
    subtype a514 is bit;
    subtype a515 is bit;
    subtype a516 is bit;
    subtype a517 is bit;
    subtype a518 is bit;
    subtype a519 is bit;
    subtype a520 is bit;
    subtype a521 is bit;
    subtype a522 is bit;
    subtype a523 is bit;
    subtype a524 is bit;
    subtype a525 is bit;
    subtype a526 is bit;
    subtype a527 is bit;
    subtype a528 is bit;
    subtype a529 is bit;
    subtype a530 is bit;
    subtype a531 is bit;
    subtype a532 is bit;
    subtype a533 is bit;
    subtype a534 is bit;
    subtype a535 is bit;
    subtype a536 is bit;
    subtype a537 is bit;
    subtype a538 is bit;
    subtype a539 is bit;
    subtype a540 is bit;
    subtype a541 is bit;
    subtype a542 is bit;
    subtype a543 is bit;
    subtype a544 is bit;
    subtype a545 is bit;
    subtype a546 is bit;
    subtype a547 is bit;
    subtype a548 is bit;
    subtype a549 is bit;
    subtype a550 is bit;
    subtype a551 is bit;
    subtype a552 is bit;
    subtype a553 is bit;
    subtype a554 is bit;
    subtype a555 is bit;
    subtype a556 is bit;
    subtype a557 is bit;
    subtype a558 is bit;
    subtype a559 is bit;
    subtype a560 is bit;
    subtype a561 is bit;
    subtype a562 is bit;
    subtype a563 is bit;
    subtype a564 is bit;
    subtype a565 is bit;
    subtype a566 is bit;
    subtype a567 is bit;
    subtype a568 is bit;
    subtype a569 is bit;
    subtype a570 is bit;
    subtype a571 is bit;
    subtype a572 is bit;
    subtype a573 is bit;
    subtype a574 is bit;
    subtype a575 is bit;
    subtype a576 is bit;
    subtype a577 is bit;
    subtype a578 is bit;
    subtype a579 is bit;
    subtype a580 is bit;
    subtype a581 is bit;
    subtype a582 is bit;
    subtype a583 is bit;
    subtype a584 is bit;
    subtype a585 is bit;
    subtype a586 is bit;
    subtype a587 is bit;
    subtype a588 is bit;
    subtype a589 is bit;
    subtype a590 is bit;
    subtype a591 is bit;
    subtype a592 is bit;
    subtype a593 is bit;
    subtype a594 is bit;
    subtype a595 is bit;
    subtype a596 is bit;
    subtype a597 is bit;
    subtype a598 is bit;
    subtype a599 is bit;
    subtype a600 is bit;
    subtype a601 is bit;
    subtype a602 is bit;
    subtype a603 is bit;
    subtype a604 is bit;
    subtype a605 is bit;
    subtype a606 is bit;
    subtype a607 is bit;
    subtype a608 is bit;
    subtype a609 is bit;
    subtype a610 is bit;
    subtype a611 is bit;
    subtype a612 is bit;
    subtype a613 is bit;
    subtype a614 is bit;
    subtype a615 is bit;
    subtype a616 is bit;
    subtype a617 is bit;
    subtype a618 is bit;
    subtype a619 is bit;
    subtype a620 is bit;
    subtype a621 is bit;
    subtype a622 is bit;
    subtype a623 is bit;
    subtype a624 is bit;
    subtype a625 is bit;
    subtype a626 is bit;
    subtype a627 is bit;
    subtype a628 is bit;
    subtype a629 is bit;
    subtype a630 is bit;
    subtype a631 is bit;
    subtype a632 is bit;
    subtype a633 is bit;
    subtype a634 is bit;
    subtype a635 is bit;
    subtype a636 is bit;
    subtype a637 is bit;
    subtype a638 is bit;
    subtype a639 is bit;
    subtype a640 is bit;
    subtype a641 is bit;
    subtype a642 is bit;
    subtype a643 is bit;
    subtype a644 is bit;
    subtype a645 is bit;
    subtype a646 is bit;
    subtype a647 is bit;
    subtype a648 is bit;
    subtype a649 is bit;
    subtype a650 is bit;
    subtype a651 is bit;
    subtype a652 is bit;
    subtype a653 is bit;
    subtype a654 is bit;
    subtype a655 is bit;
    subtype a656 is bit;
    subtype a657 is bit;
    subtype a658 is bit;
    subtype a659 is bit;
    subtype a660 is bit;
    subtype a661 is bit;
    subtype a662 is bit;
    subtype a663 is bit;
    subtype a664 is bit;
    subtype a665 is bit;
    subtype a666 is bit;
    subtype a667 is bit;
    subtype a668 is bit;
    subtype a669 is bit;
    subtype a670 is bit;
    subtype a671 is bit;
    subtype a672 is bit;
    subtype a673 is bit;
    subtype a674 is bit;
    subtype a675 is bit;
    subtype a676 is bit;
    subtype a677 is bit;
    subtype a678 is bit;
    subtype a679 is bit;
    subtype a680 is bit;
    subtype a681 is bit;
    subtype a682 is bit;
    subtype a683 is bit;
    subtype a684 is bit;
    subtype a685 is bit;
    subtype a686 is bit;
    subtype a687 is bit;
    subtype a688 is bit;
    subtype a689 is bit;
    subtype a690 is bit;
    subtype a691 is bit;
    subtype a692 is bit;
    subtype a693 is bit;
    subtype a694 is bit;
    subtype a695 is bit;
    subtype a696 is bit;
    subtype a697 is bit;
    subtype a698 is bit;
    subtype a699 is bit;
    subtype a700 is bit;
    subtype a701 is bit;
    subtype a702 is bit;
    subtype a703 is bit;
    subtype a704 is bit;
    subtype a705 is bit;
    subtype a706 is bit;
    subtype a707 is bit;
    subtype a708 is bit;
    subtype a709 is bit;
    subtype a710 is bit;
    subtype a711 is bit;
    subtype a712 is bit;
    subtype a713 is bit;
    subtype a714 is bit;
    subtype a715 is bit;
    subtype a716 is bit;
    subtype a717 is bit;
    subtype a718 is bit;
    subtype a719 is bit;
    subtype a720 is bit;
    subtype a721 is bit;
    subtype a722 is bit;
    subtype a723 is bit;
    subtype a724 is bit;
    subtype a725 is bit;
    subtype a726 is bit;
    subtype a727 is bit;
    subtype a728 is bit;
    subtype a729 is bit;
    subtype a730 is bit;
    subtype a731 is bit;
    subtype a732 is bit;
    subtype a733 is bit;
    subtype a734 is bit;
    subtype a735 is bit;
    subtype a736 is bit;
    subtype a737 is bit;
    subtype a738 is bit;
    subtype a739 is bit;
    subtype a740 is bit;
    subtype a741 is bit;
    subtype a742 is bit;
    subtype a743 is bit;
    subtype a744 is bit;
    subtype a745 is bit;
    subtype a746 is bit;
    subtype a747 is bit;
    subtype a748 is bit;
    subtype a749 is bit;
    subtype a750 is bit;
    subtype a751 is bit;
    subtype a752 is bit;
    subtype a753 is bit;
    subtype a754 is bit;
    subtype a755 is bit;
    subtype a756 is bit;
    subtype a757 is bit;
    subtype a758 is bit;
    subtype a759 is bit;
    subtype a760 is bit;
    subtype a761 is bit;
    subtype a762 is bit;
    subtype a763 is bit;
    subtype a764 is bit;
    subtype a765 is bit;
    subtype a766 is bit;
    subtype a767 is bit;
    subtype a768 is bit;
    subtype a769 is bit;
    subtype a770 is bit;
    subtype a771 is bit;
    subtype a772 is bit;
    subtype a773 is bit;
    subtype a774 is bit;
    subtype a775 is bit;
    subtype a776 is bit;
    subtype a777 is bit;
    subtype a778 is bit;
    subtype a779 is bit;
    subtype a780 is bit;
    subtype a781 is bit;
    subtype a782 is bit;
    subtype a783 is bit;
    subtype a784 is bit;
    subtype a785 is bit;
    subtype a786 is bit;
    subtype a787 is bit;
    subtype a788 is bit;
    subtype a789 is bit;
    subtype a790 is bit;
    subtype a791 is bit;
    subtype a792 is bit;
    subtype a793 is bit;
    subtype a794 is bit;
    subtype a795 is bit;
    subtype a796 is bit;
    subtype a797 is bit;
    subtype a798 is bit;
    subtype a799 is bit;
    subtype a800 is bit;
    subtype a801 is bit;
    subtype a802 is bit;
    subtype a803 is bit;
    subtype a804 is bit;
    subtype a805 is bit;
    subtype a806 is bit;
    subtype a807 is bit;
    subtype a808 is bit;
    subtype a809 is bit;
    subtype a810 is bit;
    subtype a811 is bit;
    subtype a812 is bit;
    subtype a813 is bit;
    subtype a814 is bit;
    subtype a815 is bit;
    subtype a816 is bit;
    subtype a817 is bit;
    subtype a818 is bit;
    subtype a819 is bit;
    subtype a820 is bit;
    subtype a821 is bit;
    subtype a822 is bit;
    subtype a823 is bit;
    subtype a824 is bit;
    subtype a825 is bit;
    subtype a826 is bit;
    subtype a827 is bit;
    subtype a828 is bit;
    subtype a829 is bit;
    subtype a830 is bit;
    subtype a831 is bit;
    subtype a832 is bit;
    subtype a833 is bit;
    subtype a834 is bit;
    subtype a835 is bit;
    subtype a836 is bit;
    subtype a837 is bit;
    subtype a838 is bit;
    subtype a839 is bit;
    subtype a840 is bit;
    subtype a841 is bit;
    subtype a842 is bit;
    subtype a843 is bit;
    subtype a844 is bit;
    subtype a845 is bit;
    subtype a846 is bit;
    subtype a847 is bit;
    subtype a848 is bit;
    subtype a849 is bit;
    subtype a850 is bit;
    subtype a851 is bit;
    subtype a852 is bit;
    subtype a853 is bit;
    subtype a854 is bit;
    subtype a855 is bit;
    subtype a856 is bit;
    subtype a857 is bit;
    subtype a858 is bit;
    subtype a859 is bit;
    subtype a860 is bit;
    subtype a861 is bit;
    subtype a862 is bit;
    subtype a863 is bit;
    subtype a864 is bit;
    subtype a865 is bit;
    subtype a866 is bit;
    subtype a867 is bit;
    subtype a868 is bit;
    subtype a869 is bit;
    subtype a870 is bit;
    subtype a871 is bit;
    subtype a872 is bit;
    subtype a873 is bit;
    subtype a874 is bit;
    subtype a875 is bit;
    subtype a876 is bit;
    subtype a877 is bit;
    subtype a878 is bit;
    subtype a879 is bit;
    subtype a880 is bit;
    subtype a881 is bit;
    subtype a882 is bit;
    subtype a883 is bit;
    subtype a884 is bit;
    subtype a885 is bit;
    subtype a886 is bit;
    subtype a887 is bit;
    subtype a888 is bit;
    subtype a889 is bit;
    subtype a890 is bit;
    subtype a891 is bit;
    subtype a892 is bit;
    subtype a893 is bit;
    subtype a894 is bit;
    subtype a895 is bit;
    subtype a896 is bit;
    subtype a897 is bit;
    subtype a898 is bit;
    subtype a899 is bit;
    subtype a900 is bit;
    subtype a901 is bit;
    subtype a902 is bit;
    subtype a903 is bit;
    subtype a904 is bit;
    subtype a905 is bit;
    subtype a906 is bit;
    subtype a907 is bit;
    subtype a908 is bit;
    subtype a909 is bit;
    subtype a910 is bit;
    subtype a911 is bit;
    subtype a912 is bit;
    subtype a913 is bit;
    subtype a914 is bit;
    subtype a915 is bit;
    subtype a916 is bit;
    subtype a917 is bit;
    subtype a918 is bit;
    subtype a919 is bit;
    subtype a920 is bit;
    subtype a921 is bit;
    subtype a922 is bit;
    subtype a923 is bit;
    subtype a924 is bit;
    subtype a925 is bit;
    subtype a926 is bit;
    subtype a927 is bit;
    subtype a928 is bit;
    subtype a929 is bit;
    subtype a930 is bit;
    subtype a931 is bit;
    subtype a932 is bit;
    subtype a933 is bit;
    subtype a934 is bit;
    subtype a935 is bit;
    subtype a936 is bit;
    subtype a937 is bit;
    subtype a938 is bit;
    subtype a939 is bit;
    subtype a940 is bit;
    subtype a941 is bit;
    subtype a942 is bit;
    subtype a943 is bit;
    subtype a944 is bit;
    subtype a945 is bit;
    subtype a946 is bit;
    subtype a947 is bit;
    subtype a948 is bit;
    subtype a949 is bit;
    subtype a950 is bit;
    subtype a951 is bit;
    subtype a952 is bit;
    subtype a953 is bit;
    subtype a954 is bit;
    subtype a955 is bit;
    subtype a956 is bit;
    subtype a957 is bit;
    subtype a958 is bit;
    subtype a959 is bit;
    subtype a960 is bit;
    subtype a961 is bit;
    subtype a962 is bit;
    subtype a963 is bit;
    subtype a964 is bit;
    subtype a965 is bit;
    subtype a966 is bit;
    subtype a967 is bit;
    subtype a968 is bit;
    subtype a969 is bit;
    subtype a970 is bit;
    subtype a971 is bit;
    subtype a972 is bit;
    subtype a973 is bit;
    subtype a974 is bit;
    subtype a975 is bit;
    subtype a976 is bit;
    subtype a977 is bit;
    subtype a978 is bit;
    subtype a979 is bit;
    subtype a980 is bit;
    subtype a981 is bit;
    subtype a982 is bit;
    subtype a983 is bit;
    subtype a984 is bit;
    subtype a985 is bit;
    subtype a986 is bit;
    subtype a987 is bit;
    subtype a988 is bit;
    subtype a989 is bit;
    subtype a990 is bit;
    subtype a991 is bit;
    subtype a992 is bit;
    subtype a993 is bit;
    subtype a994 is bit;
    subtype a995 is bit;
    subtype a996 is bit;
    subtype a997 is bit;
    subtype a998 is bit;
    subtype a999 is bit;
    subtype a1000 is bit;
    subtype a1001 is bit;
    subtype a1002 is bit;
    subtype a1003 is bit;
    subtype a1004 is bit;
    subtype a1005 is bit;
    subtype a1006 is bit;
    subtype a1007 is bit;
    subtype a1008 is bit;
    subtype a1009 is bit;
    subtype a1010 is bit;
    subtype a1011 is bit;
    subtype a1012 is bit;
    subtype a1013 is bit;
    subtype a1014 is bit;
    subtype a1015 is bit;
    subtype a1016 is bit;
    subtype a1017 is bit;
    subtype a1018 is bit;
    subtype a1019 is bit;
    subtype a1020 is bit;
    subtype a1021 is bit;
    subtype a1022 is bit;
    subtype a1023 is bit;
    subtype a1024 is bit;
    subtype a1025 is bit;
    subtype a1026 is bit;
    subtype a1027 is bit;
    subtype a1028 is bit;
    subtype a1029 is bit;
    subtype a1030 is bit;
    subtype a1031 is bit;
    subtype a1032 is bit;
    subtype a1033 is bit;
    subtype a1034 is bit;
    subtype a1035 is bit;
    subtype a1036 is bit;
    subtype a1037 is bit;
    subtype a1038 is bit;
    subtype a1039 is bit;
    subtype a1040 is bit;
    subtype a1041 is bit;
    subtype a1042 is bit;
    subtype a1043 is bit;
    subtype a1044 is bit;
    subtype a1045 is bit;
    subtype a1046 is bit;
    subtype a1047 is bit;
    subtype a1048 is bit;
    subtype a1049 is bit;
    subtype a1050 is bit;
    subtype a1051 is bit;
    subtype a1052 is bit;
    subtype a1053 is bit;
    subtype a1054 is bit;
    subtype a1055 is bit;
    subtype a1056 is bit;
    subtype a1057 is bit;
    subtype a1058 is bit;
    subtype a1059 is bit;
    subtype a1060 is bit;
    subtype a1061 is bit;
    subtype a1062 is bit;
    subtype a1063 is bit;
    subtype a1064 is bit;
    subtype a1065 is bit;
    subtype a1066 is bit;
    subtype a1067 is bit;
    subtype a1068 is bit;
    subtype a1069 is bit;
    subtype a1070 is bit;
    subtype a1071 is bit;
    subtype a1072 is bit;
    subtype a1073 is bit;
    subtype a1074 is bit;
    subtype a1075 is bit;
    subtype a1076 is bit;
    subtype a1077 is bit;
    subtype a1078 is bit;
    subtype a1079 is bit;
    subtype a1080 is bit;
    subtype a1081 is bit;
    subtype a1082 is bit;
    subtype a1083 is bit;
    subtype a1084 is bit;
    subtype a1085 is bit;
    subtype a1086 is bit;
    subtype a1087 is bit;
    subtype a1088 is bit;
    subtype a1089 is bit;
    subtype a1090 is bit;
    subtype a1091 is bit;
    subtype a1092 is bit;
    subtype a1093 is bit;
    subtype a1094 is bit;
    subtype a1095 is bit;
    subtype a1096 is bit;
    subtype a1097 is bit;
    subtype a1098 is bit;
    subtype a1099 is bit;
    subtype a1100 is bit;
    subtype a1101 is bit;
    subtype a1102 is bit;
    subtype a1103 is bit;
    subtype a1104 is bit;
    subtype a1105 is bit;
    subtype a1106 is bit;
    subtype a1107 is bit;
    subtype a1108 is bit;
    subtype a1109 is bit;
    subtype a1110 is bit;
    subtype a1111 is bit;
    subtype a1112 is bit;
    subtype a1113 is bit;
    subtype a1114 is bit;
    subtype a1115 is bit;
    subtype a1116 is bit;
    subtype a1117 is bit;
    subtype a1118 is bit;
    subtype a1119 is bit;
    subtype a1120 is bit;
    subtype a1121 is bit;
    subtype a1122 is bit;
    subtype a1123 is bit;
    subtype a1124 is bit;
    subtype a1125 is bit;
    subtype a1126 is bit;
    subtype a1127 is bit;
    subtype a1128 is bit;
    subtype a1129 is bit;
    subtype a1130 is bit;
    subtype a1131 is bit;
    subtype a1132 is bit;
    subtype a1133 is bit;
    subtype a1134 is bit;
    subtype a1135 is bit;
    subtype a1136 is bit;
    subtype a1137 is bit;
    subtype a1138 is bit;
    subtype a1139 is bit;
    subtype a1140 is bit;
    subtype a1141 is bit;
    subtype a1142 is bit;
    subtype a1143 is bit;
    subtype a1144 is bit;
    subtype a1145 is bit;
    subtype a1146 is bit;
    subtype a1147 is bit;
    subtype a1148 is bit;
    subtype a1149 is bit;
    subtype a1150 is bit;
    subtype a1151 is bit;
    subtype a1152 is bit;
    subtype a1153 is bit;
    subtype a1154 is bit;
    subtype a1155 is bit;
    subtype a1156 is bit;
    subtype a1157 is bit;
    subtype a1158 is bit;
    subtype a1159 is bit;
    subtype a1160 is bit;
    subtype a1161 is bit;
    subtype a1162 is bit;
    subtype a1163 is bit;
    subtype a1164 is bit;
    subtype a1165 is bit;
    subtype a1166 is bit;
    subtype a1167 is bit;
    subtype a1168 is bit;
    subtype a1169 is bit;
    subtype a1170 is bit;
    subtype a1171 is bit;
    subtype a1172 is bit;
    subtype a1173 is bit;
    subtype a1174 is bit;
    subtype a1175 is bit;
    subtype a1176 is bit;
    subtype a1177 is bit;
    subtype a1178 is bit;
    subtype a1179 is bit;
    subtype a1180 is bit;
    subtype a1181 is bit;
    subtype a1182 is bit;
    subtype a1183 is bit;
    subtype a1184 is bit;
    subtype a1185 is bit;
    subtype a1186 is bit;
    subtype a1187 is bit;
    subtype a1188 is bit;
    subtype a1189 is bit;
    subtype a1190 is bit;
    subtype a1191 is bit;
    subtype a1192 is bit;
    subtype a1193 is bit;
    subtype a1194 is bit;
    subtype a1195 is bit;
    subtype a1196 is bit;
    subtype a1197 is bit;
    subtype a1198 is bit;
    subtype a1199 is bit;
    subtype a1200 is bit;
    subtype a1201 is bit;
    subtype a1202 is bit;
    subtype a1203 is bit;
    subtype a1204 is bit;
    subtype a1205 is bit;
    subtype a1206 is bit;
    subtype a1207 is bit;
    subtype a1208 is bit;
    subtype a1209 is bit;
    subtype a1210 is bit;
    subtype a1211 is bit;
    subtype a1212 is bit;
    subtype a1213 is bit;
    subtype a1214 is bit;
    subtype a1215 is bit;
    subtype a1216 is bit;
    subtype a1217 is bit;
    subtype a1218 is bit;
    subtype a1219 is bit;
    subtype a1220 is bit;
    subtype a1221 is bit;
    subtype a1222 is bit;
    subtype a1223 is bit;
    subtype a1224 is bit;
    subtype a1225 is bit;
    subtype a1226 is bit;
    subtype a1227 is bit;
    subtype a1228 is bit;
    subtype a1229 is bit;
    subtype a1230 is bit;
    subtype a1231 is bit;
    subtype a1232 is bit;
    subtype a1233 is bit;
    subtype a1234 is bit;
    subtype a1235 is bit;
    subtype a1236 is bit;
    subtype a1237 is bit;
    subtype a1238 is bit;
    subtype a1239 is bit;
    subtype a1240 is bit;
    subtype a1241 is bit;
    subtype a1242 is bit;
    subtype a1243 is bit;
    subtype a1244 is bit;
    subtype a1245 is bit;
    subtype a1246 is bit;
    subtype a1247 is bit;
    subtype a1248 is bit;
    subtype a1249 is bit;
    subtype a1250 is bit;
    subtype a1251 is bit;
    subtype a1252 is bit;
    subtype a1253 is bit;
    subtype a1254 is bit;
    subtype a1255 is bit;
    subtype a1256 is bit;
    subtype a1257 is bit;
    subtype a1258 is bit;
    subtype a1259 is bit;
    subtype a1260 is bit;
    subtype a1261 is bit;
    subtype a1262 is bit;
    subtype a1263 is bit;
    subtype a1264 is bit;
    subtype a1265 is bit;
    subtype a1266 is bit;
    subtype a1267 is bit;
    subtype a1268 is bit;
    subtype a1269 is bit;
    subtype a1270 is bit;
    subtype a1271 is bit;
    subtype a1272 is bit;
    subtype a1273 is bit;
    subtype a1274 is bit;
    subtype a1275 is bit;
    subtype a1276 is bit;
    subtype a1277 is bit;
    subtype a1278 is bit;
    subtype a1279 is bit;
    subtype a1280 is bit;
    subtype a1281 is bit;
    subtype a1282 is bit;
    subtype a1283 is bit;
    subtype a1284 is bit;
    subtype a1285 is bit;
    subtype a1286 is bit;
    subtype a1287 is bit;
    subtype a1288 is bit;
    subtype a1289 is bit;
    subtype a1290 is bit;
    subtype a1291 is bit;
    subtype a1292 is bit;
    subtype a1293 is bit;
    subtype a1294 is bit;
    subtype a1295 is bit;
    subtype a1296 is bit;
    subtype a1297 is bit;
    subtype a1298 is bit;
    subtype a1299 is bit;
    subtype a1300 is bit;
    subtype a1301 is bit;
    subtype a1302 is bit;
    subtype a1303 is bit;
    subtype a1304 is bit;
    subtype a1305 is bit;
    subtype a1306 is bit;
    subtype a1307 is bit;
    subtype a1308 is bit;
    subtype a1309 is bit;
    subtype a1310 is bit;
    subtype a1311 is bit;
    subtype a1312 is bit;
    subtype a1313 is bit;
    subtype a1314 is bit;
    subtype a1315 is bit;
    subtype a1316 is bit;
    subtype a1317 is bit;
    subtype a1318 is bit;
    subtype a1319 is bit;
    subtype a1320 is bit;
    subtype a1321 is bit;
    subtype a1322 is bit;
    subtype a1323 is bit;
    subtype a1324 is bit;
    subtype a1325 is bit;
    subtype a1326 is bit;
    subtype a1327 is bit;
    subtype a1328 is bit;
    subtype a1329 is bit;
    subtype a1330 is bit;
    subtype a1331 is bit;
    subtype a1332 is bit;
    subtype a1333 is bit;
    subtype a1334 is bit;
    subtype a1335 is bit;
    subtype a1336 is bit;
    subtype a1337 is bit;
    subtype a1338 is bit;
    subtype a1339 is bit;
    subtype a1340 is bit;
    subtype a1341 is bit;
    subtype a1342 is bit;
    subtype a1343 is bit;
    subtype a1344 is bit;
    subtype a1345 is bit;
    subtype a1346 is bit;
    subtype a1347 is bit;
    subtype a1348 is bit;
    subtype a1349 is bit;
    subtype a1350 is bit;
    subtype a1351 is bit;
    subtype a1352 is bit;
    subtype a1353 is bit;
    subtype a1354 is bit;
    subtype a1355 is bit;
    subtype a1356 is bit;
    subtype a1357 is bit;
    subtype a1358 is bit;
    subtype a1359 is bit;
    subtype a1360 is bit;
    subtype a1361 is bit;
    subtype a1362 is bit;
    subtype a1363 is bit;
    subtype a1364 is bit;
    subtype a1365 is bit;
    subtype a1366 is bit;
    subtype a1367 is bit;
    subtype a1368 is bit;
    subtype a1369 is bit;
    subtype a1370 is bit;
    subtype a1371 is bit;
    subtype a1372 is bit;
    subtype a1373 is bit;
    subtype a1374 is bit;
    subtype a1375 is bit;
    subtype a1376 is bit;
    subtype a1377 is bit;
    subtype a1378 is bit;
    subtype a1379 is bit;
    subtype a1380 is bit;
    subtype a1381 is bit;
    subtype a1382 is bit;
    subtype a1383 is bit;
    subtype a1384 is bit;
    subtype a1385 is bit;
    subtype a1386 is bit;
    subtype a1387 is bit;
    subtype a1388 is bit;
    subtype a1389 is bit;
    subtype a1390 is bit;
    subtype a1391 is bit;
    subtype a1392 is bit;
    subtype a1393 is bit;
    subtype a1394 is bit;
    subtype a1395 is bit;
    subtype a1396 is bit;
    subtype a1397 is bit;
    subtype a1398 is bit;
    subtype a1399 is bit;
    subtype a1400 is bit;
    subtype a1401 is bit;
    subtype a1402 is bit;
    subtype a1403 is bit;
    subtype a1404 is bit;
    subtype a1405 is bit;
    subtype a1406 is bit;
    subtype a1407 is bit;
    subtype a1408 is bit;
    subtype a1409 is bit;
    subtype a1410 is bit;
    subtype a1411 is bit;
    subtype a1412 is bit;
    subtype a1413 is bit;
    subtype a1414 is bit;
    subtype a1415 is bit;
    subtype a1416 is bit;
    subtype a1417 is bit;
    subtype a1418 is bit;
    subtype a1419 is bit;
    subtype a1420 is bit;
    subtype a1421 is bit;
    subtype a1422 is bit;
    subtype a1423 is bit;
    subtype a1424 is bit;
    subtype a1425 is bit;
    subtype a1426 is bit;
    subtype a1427 is bit;
    subtype a1428 is bit;
    subtype a1429 is bit;
    subtype a1430 is bit;
    subtype a1431 is bit;
    subtype a1432 is bit;
    subtype a1433 is bit;
    subtype a1434 is bit;
    subtype a1435 is bit;
    subtype a1436 is bit;
    subtype a1437 is bit;
    subtype a1438 is bit;
    subtype a1439 is bit;
    subtype a1440 is bit;
    subtype a1441 is bit;
    subtype a1442 is bit;
    subtype a1443 is bit;
    subtype a1444 is bit;
    subtype a1445 is bit;
    subtype a1446 is bit;
    subtype a1447 is bit;
    subtype a1448 is bit;
    subtype a1449 is bit;
    subtype a1450 is bit;
    subtype a1451 is bit;
    subtype a1452 is bit;
    subtype a1453 is bit;
    subtype a1454 is bit;
    subtype a1455 is bit;
    subtype a1456 is bit;
    subtype a1457 is bit;
    subtype a1458 is bit;
    subtype a1459 is bit;
    subtype a1460 is bit;
    subtype a1461 is bit;
    subtype a1462 is bit;
    subtype a1463 is bit;
    subtype a1464 is bit;
    subtype a1465 is bit;
    subtype a1466 is bit;
    subtype a1467 is bit;
    subtype a1468 is bit;
    subtype a1469 is bit;
    subtype a1470 is bit;
    subtype a1471 is bit;
    subtype a1472 is bit;
    subtype a1473 is bit;
    subtype a1474 is bit;
    subtype a1475 is bit;
    subtype a1476 is bit;
    subtype a1477 is bit;
    subtype a1478 is bit;
    subtype a1479 is bit;
    subtype a1480 is bit;
    subtype a1481 is bit;
    subtype a1482 is bit;
    subtype a1483 is bit;
    subtype a1484 is bit;
    subtype a1485 is bit;
    subtype a1486 is bit;
    subtype a1487 is bit;
    subtype a1488 is bit;
    subtype a1489 is bit;
    subtype a1490 is bit;
    subtype a1491 is bit;
    subtype a1492 is bit;
    subtype a1493 is bit;
    subtype a1494 is bit;
    subtype a1495 is bit;
    subtype a1496 is bit;
    subtype a1497 is bit;
    subtype a1498 is bit;
    subtype a1499 is bit;
    subtype a1500 is bit;
    subtype a1501 is bit;
    subtype a1502 is bit;
    subtype a1503 is bit;
    subtype a1504 is bit;
    subtype a1505 is bit;
    subtype a1506 is bit;
    subtype a1507 is bit;
    subtype a1508 is bit;
    subtype a1509 is bit;
    subtype a1510 is bit;
    subtype a1511 is bit;
    subtype a1512 is bit;
    subtype a1513 is bit;
    subtype a1514 is bit;
    subtype a1515 is bit;
    subtype a1516 is bit;
    subtype a1517 is bit;
    subtype a1518 is bit;
    subtype a1519 is bit;
    subtype a1520 is bit;
    subtype a1521 is bit;
    subtype a1522 is bit;
    subtype a1523 is bit;
    subtype a1524 is bit;
    subtype a1525 is bit;
    subtype a1526 is bit;
    subtype a1527 is bit;
    subtype a1528 is bit;
    subtype a1529 is bit;
    subtype a1530 is bit;
    subtype a1531 is bit;
    subtype a1532 is bit;
    subtype a1533 is bit;
    subtype a1534 is bit;
    subtype a1535 is bit;
    subtype a1536 is bit;
    subtype a1537 is bit;
    subtype a1538 is bit;
    subtype a1539 is bit;
    subtype a1540 is bit;
    subtype a1541 is bit;
    subtype a1542 is bit;
    subtype a1543 is bit;
    subtype a1544 is bit;
    subtype a1545 is bit;
    subtype a1546 is bit;
    subtype a1547 is bit;
    subtype a1548 is bit;
    subtype a1549 is bit;
    subtype a1550 is bit;
    subtype a1551 is bit;
    subtype a1552 is bit;
    subtype a1553 is bit;
    subtype a1554 is bit;
    subtype a1555 is bit;
    subtype a1556 is bit;
    subtype a1557 is bit;
    subtype a1558 is bit;
    subtype a1559 is bit;
    subtype a1560 is bit;
    subtype a1561 is bit;
    subtype a1562 is bit;
    subtype a1563 is bit;
    subtype a1564 is bit;
    subtype a1565 is bit;
    subtype a1566 is bit;
    subtype a1567 is bit;
    subtype a1568 is bit;
    subtype a1569 is bit;
    subtype a1570 is bit;
    subtype a1571 is bit;
    subtype a1572 is bit;
    subtype a1573 is bit;
    subtype a1574 is bit;
    subtype a1575 is bit;
    subtype a1576 is bit;
    subtype a1577 is bit;
    subtype a1578 is bit;
    subtype a1579 is bit;
    subtype a1580 is bit;
    subtype a1581 is bit;
    subtype a1582 is bit;
    subtype a1583 is bit;
    subtype a1584 is bit;
    subtype a1585 is bit;
    subtype a1586 is bit;
    subtype a1587 is bit;
    subtype a1588 is bit;
    subtype a1589 is bit;
    subtype a1590 is bit;
    subtype a1591 is bit;
    subtype a1592 is bit;
    subtype a1593 is bit;
    subtype a1594 is bit;
    subtype a1595 is bit;
    subtype a1596 is bit;
    subtype a1597 is bit;
    subtype a1598 is bit;
    subtype a1599 is bit;
    subtype a1600 is bit;
    subtype a1601 is bit;
    subtype a1602 is bit;
    subtype a1603 is bit;
    subtype a1604 is bit;
    subtype a1605 is bit;
    subtype a1606 is bit;
    subtype a1607 is bit;
    subtype a1608 is bit;
    subtype a1609 is bit;
    subtype a1610 is bit;
    subtype a1611 is bit;
    subtype a1612 is bit;
    subtype a1613 is bit;
    subtype a1614 is bit;
    subtype a1615 is bit;
    subtype a1616 is bit;
    subtype a1617 is bit;
    subtype a1618 is bit;
    subtype a1619 is bit;
    subtype a1620 is bit;
    subtype a1621 is bit;
    subtype a1622 is bit;
    subtype a1623 is bit;
    subtype a1624 is bit;
    subtype a1625 is bit;
    subtype a1626 is bit;
    subtype a1627 is bit;
    subtype a1628 is bit;
    subtype a1629 is bit;
    subtype a1630 is bit;
    subtype a1631 is bit;
    subtype a1632 is bit;
    subtype a1633 is bit;
    subtype a1634 is bit;
    subtype a1635 is bit;
    subtype a1636 is bit;
    subtype a1637 is bit;
    subtype a1638 is bit;
    subtype a1639 is bit;
    subtype a1640 is bit;
    subtype a1641 is bit;
    subtype a1642 is bit;
    subtype a1643 is bit;
    subtype a1644 is bit;
    subtype a1645 is bit;
    subtype a1646 is bit;
    subtype a1647 is bit;
    subtype a1648 is bit;
    subtype a1649 is bit;
    subtype a1650 is bit;
    subtype a1651 is bit;
    subtype a1652 is bit;
    subtype a1653 is bit;
    subtype a1654 is bit;
    subtype a1655 is bit;
    subtype a1656 is bit;
    subtype a1657 is bit;
    subtype a1658 is bit;
    subtype a1659 is bit;
    subtype a1660 is bit;
    subtype a1661 is bit;
    subtype a1662 is bit;
    subtype a1663 is bit;
    subtype a1664 is bit;
    subtype a1665 is bit;
    subtype a1666 is bit;
    subtype a1667 is bit;
    subtype a1668 is bit;
    subtype a1669 is bit;
    subtype a1670 is bit;
    subtype a1671 is bit;
    subtype a1672 is bit;
    subtype a1673 is bit;
    subtype a1674 is bit;
    subtype a1675 is bit;
    subtype a1676 is bit;
    subtype a1677 is bit;
    subtype a1678 is bit;
    subtype a1679 is bit;
    subtype a1680 is bit;
    subtype a1681 is bit;
    subtype a1682 is bit;
    subtype a1683 is bit;
    subtype a1684 is bit;
    subtype a1685 is bit;
    subtype a1686 is bit;
    subtype a1687 is bit;
    subtype a1688 is bit;
    subtype a1689 is bit;
    subtype a1690 is bit;
    subtype a1691 is bit;
    subtype a1692 is bit;
    subtype a1693 is bit;
    subtype a1694 is bit;
    subtype a1695 is bit;
    subtype a1696 is bit;
    subtype a1697 is bit;
    subtype a1698 is bit;
    subtype a1699 is bit;
    subtype a1700 is bit;
    subtype a1701 is bit;
    subtype a1702 is bit;
    subtype a1703 is bit;
    subtype a1704 is bit;
    subtype a1705 is bit;
    subtype a1706 is bit;
    subtype a1707 is bit;
    subtype a1708 is bit;
    subtype a1709 is bit;
    subtype a1710 is bit;
    subtype a1711 is bit;
    subtype a1712 is bit;
    subtype a1713 is bit;
    subtype a1714 is bit;
    subtype a1715 is bit;
    subtype a1716 is bit;
    subtype a1717 is bit;
    subtype a1718 is bit;
    subtype a1719 is bit;
    subtype a1720 is bit;
    subtype a1721 is bit;
    subtype a1722 is bit;
    subtype a1723 is bit;
    subtype a1724 is bit;
    subtype a1725 is bit;
    subtype a1726 is bit;
    subtype a1727 is bit;
    subtype a1728 is bit;
    subtype a1729 is bit;
    subtype a1730 is bit;
    subtype a1731 is bit;
    subtype a1732 is bit;
    subtype a1733 is bit;
    subtype a1734 is bit;
    subtype a1735 is bit;
    subtype a1736 is bit;
    subtype a1737 is bit;
    subtype a1738 is bit;
    subtype a1739 is bit;
    subtype a1740 is bit;
    subtype a1741 is bit;
    subtype a1742 is bit;
    subtype a1743 is bit;
    subtype a1744 is bit;
    subtype a1745 is bit;
    subtype a1746 is bit;
    subtype a1747 is bit;
    subtype a1748 is bit;
    subtype a1749 is bit;
    subtype a1750 is bit;
    subtype a1751 is bit;
    subtype a1752 is bit;
    subtype a1753 is bit;
    subtype a1754 is bit;
    subtype a1755 is bit;
    subtype a1756 is bit;
    subtype a1757 is bit;
    subtype a1758 is bit;
    subtype a1759 is bit;
    subtype a1760 is bit;
    subtype a1761 is bit;
    subtype a1762 is bit;
    subtype a1763 is bit;
    subtype a1764 is bit;
    subtype a1765 is bit;
    subtype a1766 is bit;
    subtype a1767 is bit;
    subtype a1768 is bit;
    subtype a1769 is bit;
    subtype a1770 is bit;
    subtype a1771 is bit;
    subtype a1772 is bit;
    subtype a1773 is bit;
    subtype a1774 is bit;
    subtype a1775 is bit;
    subtype a1776 is bit;
    subtype a1777 is bit;
    subtype a1778 is bit;
    subtype a1779 is bit;
    subtype a1780 is bit;
    subtype a1781 is bit;
    subtype a1782 is bit;
    subtype a1783 is bit;
    subtype a1784 is bit;
    subtype a1785 is bit;
    subtype a1786 is bit;
    subtype a1787 is bit;
    subtype a1788 is bit;
    subtype a1789 is bit;
    subtype a1790 is bit;
    subtype a1791 is bit;
    subtype a1792 is bit;
    subtype a1793 is bit;
    subtype a1794 is bit;
    subtype a1795 is bit;
    subtype a1796 is bit;
    subtype a1797 is bit;
    subtype a1798 is bit;
    subtype a1799 is bit;
    subtype a1800 is bit;
    subtype a1801 is bit;
    subtype a1802 is bit;
    subtype a1803 is bit;
    subtype a1804 is bit;
    subtype a1805 is bit;
    subtype a1806 is bit;
    subtype a1807 is bit;
    subtype a1808 is bit;
    subtype a1809 is bit;
    subtype a1810 is bit;
    subtype a1811 is bit;
    subtype a1812 is bit;
    subtype a1813 is bit;
    subtype a1814 is bit;
    subtype a1815 is bit;
    subtype a1816 is bit;
    subtype a1817 is bit;
    subtype a1818 is bit;
    subtype a1819 is bit;
    subtype a1820 is bit;
    subtype a1821 is bit;
    subtype a1822 is bit;
    subtype a1823 is bit;
    subtype a1824 is bit;
    subtype a1825 is bit;
    subtype a1826 is bit;
    subtype a1827 is bit;
    subtype a1828 is bit;
    subtype a1829 is bit;
    subtype a1830 is bit;
    subtype a1831 is bit;
    subtype a1832 is bit;
    subtype a1833 is bit;
    subtype a1834 is bit;
    subtype a1835 is bit;
    subtype a1836 is bit;
    subtype a1837 is bit;
    subtype a1838 is bit;
    subtype a1839 is bit;
    subtype a1840 is bit;
    subtype a1841 is bit;
    subtype a1842 is bit;
    subtype a1843 is bit;
    subtype a1844 is bit;
    subtype a1845 is bit;
    subtype a1846 is bit;
    subtype a1847 is bit;
    subtype a1848 is bit;
    subtype a1849 is bit;
    subtype a1850 is bit;
    subtype a1851 is bit;
    subtype a1852 is bit;
    subtype a1853 is bit;
    subtype a1854 is bit;
    subtype a1855 is bit;
    subtype a1856 is bit;
    subtype a1857 is bit;
    subtype a1858 is bit;
    subtype a1859 is bit;
    subtype a1860 is bit;
    subtype a1861 is bit;
    subtype a1862 is bit;
    subtype a1863 is bit;
    subtype a1864 is bit;
    subtype a1865 is bit;
    subtype a1866 is bit;
    subtype a1867 is bit;
    subtype a1868 is bit;
    subtype a1869 is bit;
    subtype a1870 is bit;
    subtype a1871 is bit;
    subtype a1872 is bit;
    subtype a1873 is bit;
    subtype a1874 is bit;
    subtype a1875 is bit;
    subtype a1876 is bit;
    subtype a1877 is bit;
    subtype a1878 is bit;
    subtype a1879 is bit;
    subtype a1880 is bit;
    subtype a1881 is bit;
    subtype a1882 is bit;
    subtype a1883 is bit;
    subtype a1884 is bit;
    subtype a1885 is bit;
    subtype a1886 is bit;
    subtype a1887 is bit;
    subtype a1888 is bit;
    subtype a1889 is bit;
    subtype a1890 is bit;
    subtype a1891 is bit;
    subtype a1892 is bit;
    subtype a1893 is bit;
    subtype a1894 is bit;
    subtype a1895 is bit;
    subtype a1896 is bit;
    subtype a1897 is bit;
    subtype a1898 is bit;
    subtype a1899 is bit;
    subtype a1900 is bit;
    subtype a1901 is bit;
    subtype a1902 is bit;
    subtype a1903 is bit;
    subtype a1904 is bit;
    subtype a1905 is bit;
    subtype a1906 is bit;
    subtype a1907 is bit;
    subtype a1908 is bit;
    subtype a1909 is bit;
    subtype a1910 is bit;
    subtype a1911 is bit;
    subtype a1912 is bit;
    subtype a1913 is bit;
    subtype a1914 is bit;
    subtype a1915 is bit;
    subtype a1916 is bit;
    subtype a1917 is bit;
    subtype a1918 is bit;
    subtype a1919 is bit;
    subtype a1920 is bit;
    subtype a1921 is bit;
    subtype a1922 is bit;
    subtype a1923 is bit;
    subtype a1924 is bit;
    subtype a1925 is bit;
    subtype a1926 is bit;
    subtype a1927 is bit;
    subtype a1928 is bit;
    subtype a1929 is bit;
    subtype a1930 is bit;
    subtype a1931 is bit;
    subtype a1932 is bit;
    subtype a1933 is bit;
    subtype a1934 is bit;
    subtype a1935 is bit;
    subtype a1936 is bit;
    subtype a1937 is bit;
    subtype a1938 is bit;
    subtype a1939 is bit;
    subtype a1940 is bit;
    subtype a1941 is bit;
    subtype a1942 is bit;
    subtype a1943 is bit;
    subtype a1944 is bit;
    subtype a1945 is bit;
    subtype a1946 is bit;
    subtype a1947 is bit;
    subtype a1948 is bit;
    subtype a1949 is bit;
    subtype a1950 is bit;
    subtype a1951 is bit;
    subtype a1952 is bit;
    subtype a1953 is bit;
    subtype a1954 is bit;
    subtype a1955 is bit;
    subtype a1956 is bit;
    subtype a1957 is bit;
    subtype a1958 is bit;
    subtype a1959 is bit;
    subtype a1960 is bit;
    subtype a1961 is bit;
    subtype a1962 is bit;
    subtype a1963 is bit;
    subtype a1964 is bit;
    subtype a1965 is bit;
    subtype a1966 is bit;
    subtype a1967 is bit;
    subtype a1968 is bit;
    subtype a1969 is bit;
    subtype a1970 is bit;
    subtype a1971 is bit;
    subtype a1972 is bit;
    subtype a1973 is bit;
    subtype a1974 is bit;
    subtype a1975 is bit;
    subtype a1976 is bit;
    subtype a1977 is bit;
    subtype a1978 is bit;
    subtype a1979 is bit;
    subtype a1980 is bit;
    subtype a1981 is bit;
    subtype a1982 is bit;
    subtype a1983 is bit;
    subtype a1984 is bit;
    subtype a1985 is bit;
    subtype a1986 is bit;
    subtype a1987 is bit;
    subtype a1988 is bit;
    subtype a1989 is bit;
    subtype a1990 is bit;
    subtype a1991 is bit;
    subtype a1992 is bit;
    subtype a1993 is bit;
    subtype a1994 is bit;
    subtype a1995 is bit;
    subtype a1996 is bit;
    subtype a1997 is bit;
    subtype a1998 is bit;
    subtype a1999 is bit;
    subtype a2000 is bit;
    subtype a2001 is bit;
    subtype a2002 is bit;
    subtype a2003 is bit;
    subtype a2004 is bit;
    subtype a2005 is bit;
    subtype a2006 is bit;
    subtype a2007 is bit;
    subtype a2008 is bit;
    subtype a2009 is bit;
    subtype a2010 is bit;
    subtype a2011 is bit;
    subtype a2012 is bit;
    subtype a2013 is bit;
    subtype a2014 is bit;
    subtype a2015 is bit;
    subtype a2016 is bit;
    subtype a2017 is bit;
    subtype a2018 is bit;
    subtype a2019 is bit;
    subtype a2020 is bit;
    subtype a2021 is bit;
    subtype a2022 is bit;
    subtype a2023 is bit;
    subtype a2024 is bit;
    subtype a2025 is bit;
    subtype a2026 is bit;
    subtype a2027 is bit;
    subtype a2028 is bit;
    subtype a2029 is bit;
    subtype a2030 is bit;
    subtype a2031 is bit;
    subtype a2032 is bit;
    subtype a2033 is bit;
    subtype a2034 is bit;
    subtype a2035 is bit;
    subtype a2036 is bit;
    subtype a2037 is bit;
    subtype a2038 is bit;
    subtype a2039 is bit;
    subtype a2040 is bit;
    subtype a2041 is bit;
    subtype a2042 is bit;
    subtype a2043 is bit;
    subtype a2044 is bit;
    subtype a2045 is bit;
    subtype a2046 is bit;
    subtype a2047 is bit;
    subtype a2048 is bit;
    subtype a2049 is bit;
    subtype a2050 is bit;
    subtype a2051 is bit;
    subtype a2052 is bit;
    subtype a2053 is bit;
    subtype a2054 is bit;
    subtype a2055 is bit;
    subtype a2056 is bit;
    subtype a2057 is bit;
    subtype a2058 is bit;
    subtype a2059 is bit;
    subtype a2060 is bit;
    subtype a2061 is bit;
    subtype a2062 is bit;
    subtype a2063 is bit;
    subtype a2064 is bit;
    subtype a2065 is bit;
    subtype a2066 is bit;
    subtype a2067 is bit;
    subtype a2068 is bit;
    subtype a2069 is bit;
    subtype a2070 is bit;
    subtype a2071 is bit;
    subtype a2072 is bit;
    subtype a2073 is bit;
    subtype a2074 is bit;
    subtype a2075 is bit;
    subtype a2076 is bit;
    subtype a2077 is bit;
    subtype a2078 is bit;
    subtype a2079 is bit;
    subtype a2080 is bit;
    subtype a2081 is bit;
    subtype a2082 is bit;
    subtype a2083 is bit;
    subtype a2084 is bit;
    subtype a2085 is bit;
    subtype a2086 is bit;
    subtype a2087 is bit;
    subtype a2088 is bit;
    subtype a2089 is bit;
    subtype a2090 is bit;
    subtype a2091 is bit;
    subtype a2092 is bit;
    subtype a2093 is bit;
    subtype a2094 is bit;
    subtype a2095 is bit;
    subtype a2096 is bit;
    subtype a2097 is bit;
    subtype a2098 is bit;
    subtype a2099 is bit;
    subtype a2100 is bit;
    subtype a2101 is bit;
    subtype a2102 is bit;
    subtype a2103 is bit;
    subtype a2104 is bit;
    subtype a2105 is bit;
    subtype a2106 is bit;
    subtype a2107 is bit;
    subtype a2108 is bit;
    subtype a2109 is bit;
    subtype a2110 is bit;
    subtype a2111 is bit;
    subtype a2112 is bit;
    subtype a2113 is bit;
    subtype a2114 is bit;
    subtype a2115 is bit;
    subtype a2116 is bit;
    subtype a2117 is bit;
    subtype a2118 is bit;
    subtype a2119 is bit;
    subtype a2120 is bit;
    subtype a2121 is bit;
    subtype a2122 is bit;
    subtype a2123 is bit;
    subtype a2124 is bit;
    subtype a2125 is bit;
    subtype a2126 is bit;
    subtype a2127 is bit;
    subtype a2128 is bit;
    subtype a2129 is bit;
    subtype a2130 is bit;
    subtype a2131 is bit;
    subtype a2132 is bit;
    subtype a2133 is bit;
    subtype a2134 is bit;
    subtype a2135 is bit;
    subtype a2136 is bit;
    subtype a2137 is bit;
    subtype a2138 is bit;
    subtype a2139 is bit;
    subtype a2140 is bit;
    subtype a2141 is bit;
    subtype a2142 is bit;
    subtype a2143 is bit;
    subtype a2144 is bit;
    subtype a2145 is bit;
    subtype a2146 is bit;
    subtype a2147 is bit;
    subtype a2148 is bit;
    subtype a2149 is bit;
    subtype a2150 is bit;
    subtype a2151 is bit;
    subtype a2152 is bit;
    subtype a2153 is bit;
    subtype a2154 is bit;
    subtype a2155 is bit;
    subtype a2156 is bit;
    subtype a2157 is bit;
    subtype a2158 is bit;
    subtype a2159 is bit;
    subtype a2160 is bit;
    subtype a2161 is bit;
    subtype a2162 is bit;
    subtype a2163 is bit;
    subtype a2164 is bit;
    subtype a2165 is bit;
    subtype a2166 is bit;
    subtype a2167 is bit;
    subtype a2168 is bit;
    subtype a2169 is bit;
    subtype a2170 is bit;
    subtype a2171 is bit;
    subtype a2172 is bit;
    subtype a2173 is bit;
    subtype a2174 is bit;
    subtype a2175 is bit;
    subtype a2176 is bit;
    subtype a2177 is bit;
    subtype a2178 is bit;
    subtype a2179 is bit;
    subtype a2180 is bit;
    subtype a2181 is bit;
    subtype a2182 is bit;
    subtype a2183 is bit;
    subtype a2184 is bit;
    subtype a2185 is bit;
    subtype a2186 is bit;
    subtype a2187 is bit;
    subtype a2188 is bit;
    subtype a2189 is bit;
    subtype a2190 is bit;
    subtype a2191 is bit;
    subtype a2192 is bit;
    subtype a2193 is bit;
    subtype a2194 is bit;
    subtype a2195 is bit;
    subtype a2196 is bit;
    subtype a2197 is bit;
    subtype a2198 is bit;
    subtype a2199 is bit;
    subtype a2200 is bit;
    subtype a2201 is bit;
    subtype a2202 is bit;
    subtype a2203 is bit;
    subtype a2204 is bit;
    subtype a2205 is bit;
    subtype a2206 is bit;
    subtype a2207 is bit;
    subtype a2208 is bit;
    subtype a2209 is bit;
    subtype a2210 is bit;
    subtype a2211 is bit;
    subtype a2212 is bit;
    subtype a2213 is bit;
    subtype a2214 is bit;
    subtype a2215 is bit;
    subtype a2216 is bit;
    subtype a2217 is bit;
    subtype a2218 is bit;
    subtype a2219 is bit;
    subtype a2220 is bit;
    subtype a2221 is bit;
    subtype a2222 is bit;
    subtype a2223 is bit;
    subtype a2224 is bit;
    subtype a2225 is bit;
    subtype a2226 is bit;
    subtype a2227 is bit;
    subtype a2228 is bit;
    subtype a2229 is bit;
    subtype a2230 is bit;
    subtype a2231 is bit;
    subtype a2232 is bit;
    subtype a2233 is bit;
    subtype a2234 is bit;
    subtype a2235 is bit;
    subtype a2236 is bit;
    subtype a2237 is bit;
    subtype a2238 is bit;
    subtype a2239 is bit;
    subtype a2240 is bit;
    subtype a2241 is bit;
    subtype a2242 is bit;
    subtype a2243 is bit;
    subtype a2244 is bit;
    subtype a2245 is bit;
    subtype a2246 is bit;
    subtype a2247 is bit;
    subtype a2248 is bit;
    subtype a2249 is bit;
    subtype a2250 is bit;
    subtype a2251 is bit;
    subtype a2252 is bit;
    subtype a2253 is bit;
    subtype a2254 is bit;
    subtype a2255 is bit;
    subtype a2256 is bit;
    subtype a2257 is bit;
    subtype a2258 is bit;
    subtype a2259 is bit;
    subtype a2260 is bit;
    subtype a2261 is bit;
    subtype a2262 is bit;
    subtype a2263 is bit;
    subtype a2264 is bit;
    subtype a2265 is bit;
    subtype a2266 is bit;
    subtype a2267 is bit;
    subtype a2268 is bit;
    subtype a2269 is bit;
    subtype a2270 is bit;
    subtype a2271 is bit;
    subtype a2272 is bit;
    subtype a2273 is bit;
    subtype a2274 is bit;
    subtype a2275 is bit;
    subtype a2276 is bit;
    subtype a2277 is bit;
    subtype a2278 is bit;
    subtype a2279 is bit;
    subtype a2280 is bit;
    subtype a2281 is bit;
    subtype a2282 is bit;
    subtype a2283 is bit;
    subtype a2284 is bit;
    subtype a2285 is bit;
    subtype a2286 is bit;
    subtype a2287 is bit;
    subtype a2288 is bit;
    subtype a2289 is bit;
    subtype a2290 is bit;
    subtype a2291 is bit;
    subtype a2292 is bit;
    subtype a2293 is bit;
    subtype a2294 is bit;
    subtype a2295 is bit;
    subtype a2296 is bit;
    subtype a2297 is bit;
    subtype a2298 is bit;
    subtype a2299 is bit;
    subtype a2300 is bit;
    subtype a2301 is bit;
    subtype a2302 is bit;
    subtype a2303 is bit;
    subtype a2304 is bit;
    subtype a2305 is bit;
    subtype a2306 is bit;
    subtype a2307 is bit;
    subtype a2308 is bit;
    subtype a2309 is bit;
    subtype a2310 is bit;
    subtype a2311 is bit;
    subtype a2312 is bit;
    subtype a2313 is bit;
    subtype a2314 is bit;
    subtype a2315 is bit;
    subtype a2316 is bit;
    subtype a2317 is bit;
    subtype a2318 is bit;
    subtype a2319 is bit;
    subtype a2320 is bit;
    subtype a2321 is bit;
    subtype a2322 is bit;
    subtype a2323 is bit;
    subtype a2324 is bit;
    subtype a2325 is bit;
    subtype a2326 is bit;
    subtype a2327 is bit;
    subtype a2328 is bit;
    subtype a2329 is bit;
    subtype a2330 is bit;
    subtype a2331 is bit;
    subtype a2332 is bit;
    subtype a2333 is bit;
    subtype a2334 is bit;
    subtype a2335 is bit;
    subtype a2336 is bit;
    subtype a2337 is bit;
    subtype a2338 is bit;
    subtype a2339 is bit;
    subtype a2340 is bit;
    subtype a2341 is bit;
    subtype a2342 is bit;
    subtype a2343 is bit;
    subtype a2344 is bit;
    subtype a2345 is bit;
    subtype a2346 is bit;
    subtype a2347 is bit;
    subtype a2348 is bit;
    subtype a2349 is bit;
    subtype a2350 is bit;
    subtype a2351 is bit;
    subtype a2352 is bit;
    subtype a2353 is bit;
    subtype a2354 is bit;
    subtype a2355 is bit;
    subtype a2356 is bit;
    subtype a2357 is bit;
    subtype a2358 is bit;
    subtype a2359 is bit;
    subtype a2360 is bit;
    subtype a2361 is bit;
    subtype a2362 is bit;
    subtype a2363 is bit;
    subtype a2364 is bit;
    subtype a2365 is bit;
    subtype a2366 is bit;
    subtype a2367 is bit;
    subtype a2368 is bit;
    subtype a2369 is bit;
    subtype a2370 is bit;
    subtype a2371 is bit;
    subtype a2372 is bit;
    subtype a2373 is bit;
    subtype a2374 is bit;
    subtype a2375 is bit;
    subtype a2376 is bit;
    subtype a2377 is bit;
    subtype a2378 is bit;
    subtype a2379 is bit;
    subtype a2380 is bit;
    subtype a2381 is bit;
    subtype a2382 is bit;
    subtype a2383 is bit;
    subtype a2384 is bit;
    subtype a2385 is bit;
    subtype a2386 is bit;
    subtype a2387 is bit;
    subtype a2388 is bit;
    subtype a2389 is bit;
    subtype a2390 is bit;
    subtype a2391 is bit;
    subtype a2392 is bit;
    subtype a2393 is bit;
    subtype a2394 is bit;
    subtype a2395 is bit;
    subtype a2396 is bit;
    subtype a2397 is bit;
    subtype a2398 is bit;
    subtype a2399 is bit;
    subtype a2400 is bit;
    subtype a2401 is bit;
    subtype a2402 is bit;
    subtype a2403 is bit;
    subtype a2404 is bit;
    subtype a2405 is bit;
    subtype a2406 is bit;
    subtype a2407 is bit;
    subtype a2408 is bit;
    subtype a2409 is bit;
    subtype a2410 is bit;
    subtype a2411 is bit;
    subtype a2412 is bit;
    subtype a2413 is bit;
    subtype a2414 is bit;
    subtype a2415 is bit;
    subtype a2416 is bit;
    subtype a2417 is bit;
    subtype a2418 is bit;
    subtype a2419 is bit;
    subtype a2420 is bit;
    subtype a2421 is bit;
    subtype a2422 is bit;
    subtype a2423 is bit;
    subtype a2424 is bit;
    subtype a2425 is bit;
    subtype a2426 is bit;
    subtype a2427 is bit;
    subtype a2428 is bit;
    subtype a2429 is bit;
    subtype a2430 is bit;
    subtype a2431 is bit;
    subtype a2432 is bit;
    subtype a2433 is bit;
    subtype a2434 is bit;
    subtype a2435 is bit;
    subtype a2436 is bit;
    subtype a2437 is bit;
    subtype a2438 is bit;
    subtype a2439 is bit;
    subtype a2440 is bit;
    subtype a2441 is bit;
    subtype a2442 is bit;
    subtype a2443 is bit;
    subtype a2444 is bit;
    subtype a2445 is bit;
    subtype a2446 is bit;
    subtype a2447 is bit;
    subtype a2448 is bit;
    subtype a2449 is bit;
    subtype a2450 is bit;
    subtype a2451 is bit;
    subtype a2452 is bit;
    subtype a2453 is bit;
    subtype a2454 is bit;
    subtype a2455 is bit;
    subtype a2456 is bit;
    subtype a2457 is bit;
    subtype a2458 is bit;
    subtype a2459 is bit;
    subtype a2460 is bit;
    subtype a2461 is bit;
    subtype a2462 is bit;
    subtype a2463 is bit;
    subtype a2464 is bit;
    subtype a2465 is bit;
    subtype a2466 is bit;
    subtype a2467 is bit;
    subtype a2468 is bit;
    subtype a2469 is bit;
    subtype a2470 is bit;
    subtype a2471 is bit;
    subtype a2472 is bit;
    subtype a2473 is bit;
    subtype a2474 is bit;
    subtype a2475 is bit;
    subtype a2476 is bit;
    subtype a2477 is bit;
    subtype a2478 is bit;
    subtype a2479 is bit;
    subtype a2480 is bit;
    subtype a2481 is bit;
    subtype a2482 is bit;
    subtype a2483 is bit;
    subtype a2484 is bit;
    subtype a2485 is bit;
    subtype a2486 is bit;
    subtype a2487 is bit;
    subtype a2488 is bit;
    subtype a2489 is bit;
    subtype a2490 is bit;
    subtype a2491 is bit;
    subtype a2492 is bit;
    subtype a2493 is bit;
    subtype a2494 is bit;
    subtype a2495 is bit;
    subtype a2496 is bit;
    subtype a2497 is bit;
    subtype a2498 is bit;
    subtype a2499 is bit;
    subtype a2500 is bit;
    subtype a2501 is bit;
    subtype a2502 is bit;
    subtype a2503 is bit;
    subtype a2504 is bit;
    subtype a2505 is bit;
    subtype a2506 is bit;
    subtype a2507 is bit;
    subtype a2508 is bit;
    subtype a2509 is bit;
    subtype a2510 is bit;
    subtype a2511 is bit;
    subtype a2512 is bit;
    subtype a2513 is bit;
    subtype a2514 is bit;
    subtype a2515 is bit;
    subtype a2516 is bit;
    subtype a2517 is bit;
    subtype a2518 is bit;
    subtype a2519 is bit;
    subtype a2520 is bit;
    subtype a2521 is bit;
    subtype a2522 is bit;
    subtype a2523 is bit;
    subtype a2524 is bit;
    subtype a2525 is bit;
    subtype a2526 is bit;
    subtype a2527 is bit;
    subtype a2528 is bit;
    subtype a2529 is bit;
    subtype a2530 is bit;
    subtype a2531 is bit;
    subtype a2532 is bit;
    subtype a2533 is bit;
    subtype a2534 is bit;
    subtype a2535 is bit;
    subtype a2536 is bit;
    subtype a2537 is bit;
    subtype a2538 is bit;
    subtype a2539 is bit;
    subtype a2540 is bit;
    subtype a2541 is bit;
    subtype a2542 is bit;
    subtype a2543 is bit;
    subtype a2544 is bit;
    subtype a2545 is bit;
    subtype a2546 is bit;
    subtype a2547 is bit;
    subtype a2548 is bit;
    subtype a2549 is bit;
    subtype a2550 is bit;
    subtype a2551 is bit;
    subtype a2552 is bit;
    subtype a2553 is bit;
    subtype a2554 is bit;
    subtype a2555 is bit;
    subtype a2556 is bit;
    subtype a2557 is bit;
    subtype a2558 is bit;
    subtype a2559 is bit;
    subtype a2560 is bit;
    subtype a2561 is bit;
    subtype a2562 is bit;
    subtype a2563 is bit;
    subtype a2564 is bit;
    subtype a2565 is bit;
    subtype a2566 is bit;
    subtype a2567 is bit;
    subtype a2568 is bit;
    subtype a2569 is bit;
    subtype a2570 is bit;
    subtype a2571 is bit;
    subtype a2572 is bit;
    subtype a2573 is bit;
    subtype a2574 is bit;
    subtype a2575 is bit;
    subtype a2576 is bit;
    subtype a2577 is bit;
    subtype a2578 is bit;
    subtype a2579 is bit;
    subtype a2580 is bit;
    subtype a2581 is bit;
    subtype a2582 is bit;
    subtype a2583 is bit;
    subtype a2584 is bit;
    subtype a2585 is bit;
    subtype a2586 is bit;
    subtype a2587 is bit;
    subtype a2588 is bit;
    subtype a2589 is bit;
    subtype a2590 is bit;
    subtype a2591 is bit;
    subtype a2592 is bit;
    subtype a2593 is bit;
    subtype a2594 is bit;
    subtype a2595 is bit;
    subtype a2596 is bit;
    subtype a2597 is bit;
    subtype a2598 is bit;
    subtype a2599 is bit;
    subtype a2600 is bit;
    subtype a2601 is bit;
    subtype a2602 is bit;
    subtype a2603 is bit;
    subtype a2604 is bit;
    subtype a2605 is bit;
    subtype a2606 is bit;
    subtype a2607 is bit;
    subtype a2608 is bit;
    subtype a2609 is bit;
    subtype a2610 is bit;
    subtype a2611 is bit;
    subtype a2612 is bit;
    subtype a2613 is bit;
    subtype a2614 is bit;
    subtype a2615 is bit;
    subtype a2616 is bit;
    subtype a2617 is bit;
    subtype a2618 is bit;
    subtype a2619 is bit;
    subtype a2620 is bit;
    subtype a2621 is bit;
    subtype a2622 is bit;
    subtype a2623 is bit;
    subtype a2624 is bit;
    subtype a2625 is bit;
    subtype a2626 is bit;
    subtype a2627 is bit;
    subtype a2628 is bit;
    subtype a2629 is bit;
    subtype a2630 is bit;
    subtype a2631 is bit;
    subtype a2632 is bit;
    subtype a2633 is bit;
    subtype a2634 is bit;
    subtype a2635 is bit;
    subtype a2636 is bit;
    subtype a2637 is bit;
    subtype a2638 is bit;
    subtype a2639 is bit;
    subtype a2640 is bit;
    subtype a2641 is bit;
    subtype a2642 is bit;
    subtype a2643 is bit;
    subtype a2644 is bit;
    subtype a2645 is bit;
    subtype a2646 is bit;
    subtype a2647 is bit;
    subtype a2648 is bit;
    subtype a2649 is bit;
    subtype a2650 is bit;
    subtype a2651 is bit;
    subtype a2652 is bit;
    subtype a2653 is bit;
    subtype a2654 is bit;
    subtype a2655 is bit;
    subtype a2656 is bit;
    subtype a2657 is bit;
    subtype a2658 is bit;
    subtype a2659 is bit;
    subtype a2660 is bit;
    subtype a2661 is bit;
    subtype a2662 is bit;
    subtype a2663 is bit;
    subtype a2664 is bit;
    subtype a2665 is bit;
    subtype a2666 is bit;
    subtype a2667 is bit;
    subtype a2668 is bit;
    subtype a2669 is bit;
    subtype a2670 is bit;
end package c;
