library ieee;use ieee.numeric_std.all;use ieee.std_logic_1164.all;entity t is generic(type s;z:boolean:=false);port(l:std'l);end;architecture a of t is type t is array(0)of t;signal r:r range 0 to 0;signal d:r range 0 to 0;signal d:n;begin y<='0'when(0)and 0 else'0';m(0);process(l)begin
if(0)then if 0 then w<=0;end if;if 0 then
r<=0;end if;end if;end process;end;