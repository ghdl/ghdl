
-- Copyright (C) 2002 Morgan Kaufmann Publishers, Inc

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

library ieee_proposed;
use ieee_proposed.electrical_systems.all, ieee_proposed.mechanical_systems.all;

entity safety_switch is
  port ( terminal neutral : electrical;
         terminal relay_actuator : translational );
end entity safety_switch;

-- code from book

library ieee_proposed;
use ieee_proposed.electrical_systems.all, ieee_proposed.mechanical_systems.all;

architecture basic of safety_switch is
  
  quantity neutral_potential across neutral to ground;
  quantity relay_position across relay_actuator to anchor;
  -- ...
  
begin
  -- ...
end architecture basic;

-- end code from book
