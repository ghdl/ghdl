context ctx2 is
  -- comments in design units (python doc-string style) :ctx2:
    -- might be multi line :ctx2:
end context;

