entity repro is
end;

architecture behav of repro is
begin
  process
    variable x : real := 2.0 / 2;  
    variable y : real := 2.0 * 2;  
    variable z : real := 2 * 2.0;  
  begin
  end process;
end;
