architecture package