package pkg is
-- function identifier return integer;
 procedure identifier;
 alias identifier_alias_fun is identifier[return integer];
-- alias identifier_alias_proc is identifier[];
end package; 
