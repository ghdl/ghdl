package--
function is if('t �';