architecture function is;0package