package
function begin if a r';