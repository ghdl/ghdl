entity e4 is end;

architecture a of e4 is
begin
    process
    begin
        report "" severity note;
    end process;
end;
