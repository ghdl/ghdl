library ieee;
use ieee.std_logic_1164.all;

entity example is
  generic (
    PARAMETER : std_logic_vector(7 downto 0));
end example;

architecture behavioral of example is
begin
end behavioral;
