use std.textio.all;

entity t1 is
end;

architecture behav of t1 is
  subtype stext is text;
begin
end behav;
