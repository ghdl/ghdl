entity ent is
end;

architecture arch of ent is
begin
end;
