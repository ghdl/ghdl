entity sig1 is
end;

use work.pkg.all;

architecture behav of sig1 is
  signal s : rec_4;
begin
end behav;
