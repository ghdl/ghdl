architecture 0for(""x""4000000000x"