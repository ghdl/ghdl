package pkg2 is
  function f (a : integer) return integer;
  function f (a : integer) return integer;
end pkg2;
