library ieee;
use ieee.std_logic_1164.all;

library ieee;
use ieee.numeric_std.all;

entity fsm_23 is
	port (
		clock : in  std_logic;
		reset : in  std_logic;
		in0 : in  std_logic;
		out181 : out std_logic;
		out182 : out std_logic;
		out183 : out std_logic;
		out184 : out std_logic;
		out185 : out std_logic;
		out8 : out std_logic;
		out13 : out std_logic;
		out14 : out std_logic;
		out16 : out std_logic;
		out18 : out std_logic;
		out19 : out std_logic;
		out20 : out std_logic;
		out21 : out std_logic;
		out22 : out std_logic;
		in2 : in  std_logic;
		out23 : out std_logic;
		out24 : out std_logic;
		out25 : out std_logic;
		out26 : out std_logic;
		out27 : out std_logic;
		out28 : out std_logic;
		out29 : out std_logic;
		out30 : out std_logic;
		out31 : out std_logic;
		out33 : out std_logic;
		out35 : out std_logic;
		out36 : out std_logic;
		out38 : out std_logic;
		out40 : out std_logic;
		out42 : out std_logic;
		in3 : in  std_logic;
		out44 : out std_logic;
		out46 : out std_logic;
		out48 : out std_logic;
		out49 : out std_logic;
		out50 : out std_logic;
		out52 : out std_logic;
		out54 : out std_logic;
		out56 : out std_logic;
		out57 : out std_logic;
		out58 : out std_logic;
		in4 : in  std_logic;
		out60 : out std_logic;
		in5 : in  std_logic;
		out164 : out std_logic;
		out165 : out std_logic;
		out167 : out std_logic;
		out168 : out std_logic;
		out170 : out std_logic;
		out171 : out std_logic;
		out173 : out std_logic;
		out174 : out std_logic;
		out176 : out std_logic;
		out178 : out std_logic;
		out0 : out std_logic;
		out1 : out std_logic;
		out2 : out std_logic;
		in1 : in  std_logic;
		out4 : out std_logic;
		out90 : out std_logic;
		out91 : out std_logic;
		out97 : out std_logic;
		out99 : out std_logic;
		out101 : out std_logic;
		in6 : in  std_logic;
		out103 : out std_logic;
		out105 : out std_logic;
		out106 : out std_logic;
		out107 : out std_logic;
		out108 : out std_logic;
		out135 : out std_logic;
		out136 : out std_logic;
		out137 : out std_logic;
		out138 : out std_logic;
		in11 : in  std_logic;
		out140 : out std_logic;
		out141 : out std_logic;
		out142 : out std_logic;
		out143 : out std_logic;
		out145 : out std_logic;
		out146 : out std_logic;
		out148 : out std_logic;
		out150 : out std_logic;
		out153 : out std_logic;
		out154 : out std_logic;
		out155 : out std_logic;
		out156 : out std_logic;
		out157 : out std_logic;
		out158 : out std_logic;
		out159 : out std_logic;
		out160 : out std_logic;
		out161 : out std_logic;
		out162 : out std_logic;
		out111 : out std_logic;
		out112 : out std_logic;
		out114 : out std_logic;
		out116 : out std_logic;
		out118 : out std_logic;
		out120 : out std_logic;
		out121 : out std_logic;
		out122 : out std_logic;
		out123 : out std_logic;
		out124 : out std_logic;
		out125 : out std_logic;
		out126 : out std_logic;
		in7 : in  std_logic;
		out129 : out std_logic;
		out130 : out std_logic;
		in8 : in  std_logic;
		out131 : out std_logic;
		in9 : in  std_logic;
		out132 : out std_logic;
		out133 : out std_logic;
		out134 : out std_logic;
		in10 : in  std_logic;
		out186 : out std_logic;
		out187 : out std_logic;
		out190 : out std_logic;
		out195 : out std_logic;
		out197 : out std_logic;
		out198 : out std_logic;
		out199 : out std_logic;
		out200 : out std_logic;
		out201 : out std_logic;
		out203 : out std_logic;
		out204 : out std_logic;
		out206 : out std_logic;
		out207 : out std_logic;
		out209 : out std_logic;
		out210 : out std_logic;
		out212 : out std_logic;
		out213 : out std_logic;
		out215 : out std_logic;
		out217 : out std_logic;
		out220 : out std_logic;
		out221 : out std_logic;
		out222 : out std_logic;
		out223 : out std_logic;
		out224 : out std_logic;
		out225 : out std_logic;
		out226 : out std_logic;
		out227 : out std_logic;
		out228 : out std_logic;
		out229 : out std_logic;
		out231 : out std_logic;
		out232 : out std_logic;
		out234 : out std_logic;
		out235 : out std_logic;
		out237 : out std_logic;
		out238 : out std_logic;
		out240 : out std_logic;
		out241 : out std_logic;
		out243 : out std_logic;
		out245 : out std_logic;
		out248 : out std_logic;
		out249 : out std_logic;
		out250 : out std_logic;
		out251 : out std_logic;
		out252 : out std_logic;
		out253 : out std_logic;
		out254 : out std_logic;
		out255 : out std_logic;
		out256 : out std_logic;
		out257 : out std_logic;
		out259 : out std_logic;
		out260 : out std_logic;
		out262 : out std_logic;
		out263 : out std_logic;
		out265 : out std_logic;
		out266 : out std_logic;
		out268 : out std_logic;
		out269 : out std_logic;
		out271 : out std_logic;
		out273 : out std_logic;
		out276 : out std_logic;
		out277 : out std_logic;
		out278 : out std_logic;
		out279 : out std_logic;
		out280 : out std_logic;
		out281 : out std_logic;
		out282 : out std_logic;
		out283 : out std_logic;
		out284 : out std_logic;
		out285 : out std_logic;
		out286 : out std_logic;
		out287 : out std_logic;
		out288 : out std_logic;
		out289 : out std_logic;
		out290 : out std_logic;
		out291 : out std_logic;
		out292 : out std_logic;
		out293 : out std_logic;
		out294 : out std_logic;
		out295 : out std_logic;
		out296 : out std_logic;
		out297 : out std_logic;
		out298 : out std_logic;
		out311 : out std_logic;
		out312 : out std_logic;
		out313 : out std_logic;
		out314 : out std_logic;
		out315 : out std_logic;
		out316 : out std_logic;
		out318 : out std_logic;
		out321 : out std_logic;
		out322 : out std_logic;
		out323 : out std_logic;
		out324 : out std_logic;
		out325 : out std_logic;
		out326 : out std_logic;
		out327 : out std_logic;
		out328 : out std_logic;
		out329 : out std_logic;
		out333 : out std_logic;
		out341 : out std_logic;
		out342 : out std_logic;
		out343 : out std_logic;
		out344 : out std_logic;
		out345 : out std_logic;
		out346 : out std_logic;
		out349 : out std_logic;
		out350 : out std_logic;
		out351 : out std_logic;
		out352 : out std_logic;
		out353 : out std_logic;
		out354 : out std_logic;
		out355 : out std_logic;
		out357 : out std_logic;
		out361 : out std_logic;
		out362 : out std_logic;
		out363 : out std_logic;
		out364 : out std_logic;
		out366 : out std_logic;
		out367 : out std_logic;
		out371 : out std_logic;
		out372 : out std_logic;
		out373 : out std_logic;
		out382 : out std_logic;
		out383 : out std_logic;
		out385 : out std_logic;
		out393 : out std_logic;
		out394 : out std_logic;
		out395 : out std_logic;
		out396 : out std_logic;
		out398 : out std_logic;
		out400 : out std_logic;
		out401 : out std_logic;
		out402 : out std_logic;
		out404 : out std_logic;
		out406 : out std_logic;
		out407 : out std_logic;
		out408 : out std_logic;
		out409 : out std_logic;
		out410 : out std_logic;
		out411 : out std_logic;
		out412 : out std_logic;
		out413 : out std_logic;
		out414 : out std_logic;
		out416 : out std_logic;
		out417 : out std_logic;
		out418 : out std_logic;
		out419 : out std_logic;
		out422 : out std_logic;
		out423 : out std_logic;
		out425 : out std_logic;
		out426 : out std_logic;
		out428 : out std_logic;
		out429 : out std_logic;
		out430 : out std_logic;
		out431 : out std_logic;
		out433 : out std_logic;
		out434 : out std_logic;
		out435 : out std_logic;
		out436 : out std_logic;
		out437 : out std_logic;
		out438 : out std_logic;
		out440 : out std_logic;
		out441 : out std_logic;
		out443 : out std_logic;
		out444 : out std_logic;
		out445 : out std_logic;
		out446 : out std_logic;
		out447 : out std_logic;
		out450 : out std_logic;
		out451 : out std_logic;
		out454 : out std_logic;
		out455 : out std_logic;
		out457 : out std_logic;
		out458 : out std_logic;
		out459 : out std_logic;
		out460 : out std_logic;
		out461 : out std_logic;
		out462 : out std_logic;
		out463 : out std_logic;
		out464 : out std_logic;
		out465 : out std_logic;
		out466 : out std_logic;
		out467 : out std_logic;
		out468 : out std_logic;
		out469 : out std_logic;
		out472 : out std_logic;
		out475 : out std_logic;
		out481 : out std_logic;
		out482 : out std_logic;
		out483 : out std_logic;
		out484 : out std_logic;
		out487 : out std_logic;
		out488 : out std_logic;
		out491 : out std_logic;
		out495 : out std_logic;
		out496 : out std_logic;
		out497 : out std_logic;
		out498 : out std_logic;
		out499 : out std_logic;
		out500 : out std_logic;
		out501 : out std_logic;
		out512 : out std_logic;
		out513 : out std_logic;
		out517 : out std_logic;
		out518 : out std_logic;
		out519 : out std_logic;
		out521 : out std_logic;
		out522 : out std_logic;
		out524 : out std_logic;
		out525 : out std_logic;
		out526 : out std_logic;
		out527 : out std_logic;
		out528 : out std_logic;
		out531 : out std_logic;
		out540 : out std_logic;
		out542 : out std_logic;
		out544 : out std_logic;
		out545 : out std_logic;
		out554 : out std_logic;
		out555 : out std_logic;
		out559 : out std_logic;
		out560 : out std_logic;
		out561 : out std_logic;
		out562 : out std_logic;
		out563 : out std_logic;
		out566 : out std_logic;
		out567 : out std_logic;
		out570 : out std_logic;
		out572 : out std_logic;
		out575 : out std_logic;
		out577 : out std_logic;
		out578 : out std_logic;
		out580 : out std_logic;
		out581 : out std_logic
	);
end fsm_23;

architecture augh of fsm_23 is

	signal state_cur  : std_logic_vector(0 to 240) := (7 => '1', others => '0');
	signal state_next : std_logic_vector(0 to 240) := (7 => '1', others => '0');

	-- Buffers for outputs
	signal out122_buf : std_logic := '0';
	signal out122_bufn : std_logic;
	signal out36_buf : std_logic := '0';
	signal out36_bufn : std_logic;
	signal out49_buf : std_logic := '0';
	signal out49_bufn : std_logic;
	signal out35_buf : std_logic := '0';
	signal out35_bufn : std_logic;
	signal out27_buf : std_logic := '0';
	signal out27_bufn : std_logic;
	signal out16_buf : std_logic := '0';
	signal out16_bufn : std_logic;
	signal out25_buf : std_logic := '0';
	signal out25_bufn : std_logic;
	signal out20_buf : std_logic := '0';
	signal out20_bufn : std_logic;
	signal out57_buf : std_logic := '0';
	signal out57_bufn : std_logic;
	signal out23_buf : std_logic := '0';
	signal out23_bufn : std_logic;
	signal out136_buf : std_logic := '0';
	signal out136_bufn : std_logic;
	signal out0_buf : std_logic := '0';
	signal out0_bufn : std_logic;
	signal out134_buf : std_logic := '0';
	signal out134_bufn : std_logic;
	signal out13_buf : std_logic := '0';
	signal out13_bufn : std_logic;
	signal out131_buf : std_logic := '0';
	signal out131_bufn : std_logic;
	signal out129_buf : std_logic := '0';
	signal out129_bufn : std_logic;
	signal out111_buf : std_logic := '0';
	signal out111_bufn : std_logic;
	signal out31_buf : std_logic := '0';
	signal out31_bufn : std_logic;
	signal out126_buf : std_logic := '0';
	signal out126_bufn : std_logic;
	signal out106_buf : std_logic := '0';
	signal out106_bufn : std_logic;
	signal out124_buf : std_logic := '0';
	signal out124_bufn : std_logic;
	signal out138_buf : std_logic := '0';
	signal out138_bufn : std_logic;
	signal out141_buf : std_logic := '0';
	signal out141_bufn : std_logic;
	signal out143_buf : std_logic := '0';
	signal out143_bufn : std_logic;
	signal out146_buf : std_logic := '0';
	signal out146_bufn : std_logic;
	signal out150_buf : std_logic := '0';
	signal out150_bufn : std_logic;
	signal out153_buf : std_logic := '0';
	signal out153_bufn : std_logic;
	signal out155_buf : std_logic := '0';
	signal out155_bufn : std_logic;
	signal out158_buf : std_logic := '0';
	signal out158_bufn : std_logic;
	signal out162_buf : std_logic := '0';
	signal out162_bufn : std_logic;
	signal out165_buf : std_logic := '0';
	signal out165_bufn : std_logic;
	signal out168_buf : std_logic := '0';
	signal out168_bufn : std_logic;
	signal out171_buf : std_logic := '0';
	signal out171_bufn : std_logic;
	signal out174_buf : std_logic := '0';
	signal out174_bufn : std_logic;
	signal out178_buf : std_logic := '0';
	signal out178_bufn : std_logic;
	signal out181_buf : std_logic := '0';
	signal out181_bufn : std_logic;
	signal out183_buf : std_logic := '0';
	signal out183_bufn : std_logic;
	signal out197_buf : std_logic := '0';
	signal out197_bufn : std_logic;
	signal out201_buf : std_logic := '0';
	signal out201_bufn : std_logic;
	signal out204_buf : std_logic := '0';
	signal out204_bufn : std_logic;
	signal out207_buf : std_logic := '0';
	signal out207_bufn : std_logic;
	signal out210_buf : std_logic := '0';
	signal out210_bufn : std_logic;
	signal out213_buf : std_logic := '0';
	signal out213_bufn : std_logic;
	signal out217_buf : std_logic := '0';
	signal out217_bufn : std_logic;
	signal out220_buf : std_logic := '0';
	signal out220_bufn : std_logic;
	signal out222_buf : std_logic := '0';
	signal out222_bufn : std_logic;
	signal out225_buf : std_logic := '0';
	signal out225_bufn : std_logic;
	signal out229_buf : std_logic := '0';
	signal out229_bufn : std_logic;
	signal out232_buf : std_logic := '0';
	signal out232_bufn : std_logic;
	signal out235_buf : std_logic := '0';
	signal out235_bufn : std_logic;
	signal out238_buf : std_logic := '0';
	signal out238_bufn : std_logic;
	signal out241_buf : std_logic := '0';
	signal out241_bufn : std_logic;
	signal out245_buf : std_logic := '0';
	signal out245_bufn : std_logic;
	signal out248_buf : std_logic := '0';
	signal out248_bufn : std_logic;
	signal out250_buf : std_logic := '0';
	signal out250_bufn : std_logic;
	signal out253_buf : std_logic := '0';
	signal out253_bufn : std_logic;
	signal out257_buf : std_logic := '0';
	signal out257_bufn : std_logic;
	signal out260_buf : std_logic := '0';
	signal out260_bufn : std_logic;
	signal out263_buf : std_logic := '0';
	signal out263_bufn : std_logic;
	signal out266_buf : std_logic := '0';
	signal out266_bufn : std_logic;
	signal out269_buf : std_logic := '0';
	signal out269_bufn : std_logic;
	signal out273_buf : std_logic := '0';
	signal out273_bufn : std_logic;
	signal out276_buf : std_logic := '0';
	signal out276_bufn : std_logic;
	signal out278_buf : std_logic := '0';
	signal out278_bufn : std_logic;
	signal out280_buf : std_logic := '0';
	signal out280_bufn : std_logic;
	signal out281_buf : std_logic := '0';
	signal out281_bufn : std_logic;
	signal out282_buf : std_logic := '0';
	signal out282_bufn : std_logic;
	signal out284_buf : std_logic := '0';
	signal out284_bufn : std_logic;
	signal out285_buf : std_logic := '0';
	signal out285_bufn : std_logic;
	signal out287_buf : std_logic := '0';
	signal out287_bufn : std_logic;
	signal out288_buf : std_logic := '0';
	signal out288_bufn : std_logic;
	signal out289_buf : std_logic := '0';
	signal out289_bufn : std_logic;
	signal out290_buf : std_logic := '0';
	signal out290_bufn : std_logic;
	signal out291_buf : std_logic := '0';
	signal out291_bufn : std_logic;
	signal out292_buf : std_logic := '0';
	signal out292_bufn : std_logic;
	signal out293_buf : std_logic := '0';
	signal out293_bufn : std_logic;
	signal out294_buf : std_logic := '0';
	signal out294_bufn : std_logic;
	signal out295_buf : std_logic := '0';
	signal out295_bufn : std_logic;
	signal out296_buf : std_logic := '0';
	signal out296_bufn : std_logic;
	signal out312_buf : std_logic := '0';
	signal out312_bufn : std_logic;
	signal out313_buf : std_logic := '0';
	signal out313_bufn : std_logic;
	signal out314_buf : std_logic := '0';
	signal out314_bufn : std_logic;
	signal out315_buf : std_logic := '0';
	signal out315_bufn : std_logic;
	signal out318_buf : std_logic := '0';
	signal out318_bufn : std_logic;
	signal out322_buf : std_logic := '0';
	signal out322_bufn : std_logic;
	signal out323_buf : std_logic := '0';
	signal out323_bufn : std_logic;
	signal out324_buf : std_logic := '0';
	signal out324_bufn : std_logic;
	signal out325_buf : std_logic := '0';
	signal out325_bufn : std_logic;
	signal out326_buf : std_logic := '0';
	signal out326_bufn : std_logic;
	signal out327_buf : std_logic := '0';
	signal out327_bufn : std_logic;
	signal out328_buf : std_logic := '0';
	signal out328_bufn : std_logic;
	signal out333_buf : std_logic := '0';
	signal out333_bufn : std_logic;
	signal out341_buf : std_logic := '0';
	signal out341_bufn : std_logic;
	signal out342_buf : std_logic := '0';
	signal out342_bufn : std_logic;
	signal out343_buf : std_logic := '0';
	signal out343_bufn : std_logic;
	signal out344_buf : std_logic := '0';
	signal out344_bufn : std_logic;
	signal out346_buf : std_logic := '0';
	signal out346_bufn : std_logic;
	signal out349_buf : std_logic := '0';
	signal out349_bufn : std_logic;
	signal out351_buf : std_logic := '0';
	signal out351_bufn : std_logic;
	signal out352_buf : std_logic := '0';
	signal out352_bufn : std_logic;
	signal out353_buf : std_logic := '0';
	signal out353_bufn : std_logic;
	signal out354_buf : std_logic := '0';
	signal out354_bufn : std_logic;
	signal out357_buf : std_logic := '0';
	signal out357_bufn : std_logic;
	signal out361_buf : std_logic := '0';
	signal out361_bufn : std_logic;
	signal out364_buf : std_logic := '0';
	signal out364_bufn : std_logic;
	signal out366_buf : std_logic := '0';
	signal out366_bufn : std_logic;
	signal out371_buf : std_logic := '0';
	signal out371_bufn : std_logic;
	signal out393_buf : std_logic := '0';
	signal out393_bufn : std_logic;
	signal out394_buf : std_logic := '0';
	signal out394_bufn : std_logic;
	signal out395_buf : std_logic := '0';
	signal out395_bufn : std_logic;
	signal out400_buf : std_logic := '0';
	signal out400_bufn : std_logic;
	signal out401_buf : std_logic := '0';
	signal out401_bufn : std_logic;
	signal out404_buf : std_logic := '0';
	signal out404_bufn : std_logic;
	signal out407_buf : std_logic := '0';
	signal out407_bufn : std_logic;
	signal out408_buf : std_logic := '0';
	signal out408_bufn : std_logic;
	signal out409_buf : std_logic := '0';
	signal out409_bufn : std_logic;
	signal out410_buf : std_logic := '0';
	signal out410_bufn : std_logic;
	signal out413_buf : std_logic := '0';
	signal out413_bufn : std_logic;
	signal out414_buf : std_logic := '0';
	signal out414_bufn : std_logic;
	signal out417_buf : std_logic := '0';
	signal out417_bufn : std_logic;
	signal out418_buf : std_logic := '0';
	signal out418_bufn : std_logic;
	signal out422_buf : std_logic := '0';
	signal out422_bufn : std_logic;
	signal out426_buf : std_logic := '0';
	signal out426_bufn : std_logic;
	signal out428_buf : std_logic := '0';
	signal out428_bufn : std_logic;
	signal out431_buf : std_logic := '0';
	signal out431_bufn : std_logic;
	signal out433_buf : std_logic := '0';
	signal out433_bufn : std_logic;
	signal out434_buf : std_logic := '0';
	signal out434_bufn : std_logic;
	signal out435_buf : std_logic := '0';
	signal out435_bufn : std_logic;
	signal out436_buf : std_logic := '0';
	signal out436_bufn : std_logic;
	signal out437_buf : std_logic := '0';
	signal out437_bufn : std_logic;
	signal out438_buf : std_logic := '0';
	signal out438_bufn : std_logic;
	signal out440_buf : std_logic := '0';
	signal out440_bufn : std_logic;
	signal out444_buf : std_logic := '0';
	signal out444_bufn : std_logic;
	signal out446_buf : std_logic := '0';
	signal out446_bufn : std_logic;
	signal out451_buf : std_logic := '0';
	signal out451_bufn : std_logic;
	signal out457_buf : std_logic := '0';
	signal out457_bufn : std_logic;
	signal out458_buf : std_logic := '0';
	signal out458_bufn : std_logic;
	signal out459_buf : std_logic := '0';
	signal out459_bufn : std_logic;
	signal out460_buf : std_logic := '0';
	signal out460_bufn : std_logic;
	signal out461_buf : std_logic := '0';
	signal out461_bufn : std_logic;
	signal out463_buf : std_logic := '0';
	signal out463_bufn : std_logic;
	signal out464_buf : std_logic := '0';
	signal out464_bufn : std_logic;
	signal out466_buf : std_logic := '0';
	signal out466_bufn : std_logic;
	signal out468_buf : std_logic := '0';
	signal out468_bufn : std_logic;
	signal out472_buf : std_logic := '0';
	signal out472_bufn : std_logic;
	signal out475_buf : std_logic := '0';
	signal out475_bufn : std_logic;
	signal out481_buf : std_logic := '0';
	signal out481_bufn : std_logic;
	signal out482_buf : std_logic := '0';
	signal out482_bufn : std_logic;
	signal out483_buf : std_logic := '0';
	signal out483_bufn : std_logic;
	signal out487_buf : std_logic := '0';
	signal out487_bufn : std_logic;
	signal out495_buf : std_logic := '0';
	signal out495_bufn : std_logic;
	signal out496_buf : std_logic := '0';
	signal out496_bufn : std_logic;
	signal out497_buf : std_logic := '0';
	signal out497_bufn : std_logic;
	signal out499_buf : std_logic := '0';
	signal out499_bufn : std_logic;
	signal out500_buf : std_logic := '0';
	signal out500_bufn : std_logic;
	signal out512_buf : std_logic := '0';
	signal out512_bufn : std_logic;
	signal out517_buf : std_logic := '0';
	signal out517_bufn : std_logic;
	signal out518_buf : std_logic := '0';
	signal out518_bufn : std_logic;
	signal out521_buf : std_logic := '0';
	signal out521_bufn : std_logic;
	signal out524_buf : std_logic := '0';
	signal out524_bufn : std_logic;
	signal out525_buf : std_logic := '0';
	signal out525_bufn : std_logic;
	signal out526_buf : std_logic := '0';
	signal out526_bufn : std_logic;
	signal out531_buf : std_logic := '0';
	signal out531_bufn : std_logic;
	signal out554_buf : std_logic := '0';
	signal out554_bufn : std_logic;
	signal out562_buf : std_logic := '0';
	signal out562_bufn : std_logic;
	signal out566_buf : std_logic := '0';
	signal out566_bufn : std_logic;

	-- Retiming: counters
	signal rtmcounter0 :      unsigned(4 downto 0) := (others => '0');
	signal rtmcounter0_next : unsigned(4 downto 0);

	-- Retiming: Output of comparators
	signal rtmcmp90 : std_logic;
	signal rtmcmp95 : std_logic;
	signal rtmcmp98 : std_logic;
	signal rtmcmp104 : std_logic;
	signal rtmcmp148 : std_logic;
	signal rtmcmp167 : std_logic;
	signal rtmcmp174 : std_logic;
	signal rtmcmp181 : std_logic;
	signal rtmcmp183 : std_logic;
	signal rtmcmp194 : std_logic;
	signal rtmcmp197 : std_logic;
	signal rtmcmp203 : std_logic;
	signal rtmcmp205 : std_logic;
	signal rtmcmp215 : std_logic;

	-- Function calls: return IDs

begin

	-- Sequential process
	-- Set the current state

	process (clock)
	begin
		if rising_edge(clock) then

			-- Next state
			state_cur <= state_next;
			-- Buffers for outputs
			out122_buf <= out122_bufn;
			out36_buf <= out36_bufn;
			out49_buf <= out49_bufn;
			out35_buf <= out35_bufn;
			out27_buf <= out27_bufn;
			out16_buf <= out16_bufn;
			out25_buf <= out25_bufn;
			out20_buf <= out20_bufn;
			out57_buf <= out57_bufn;
			out23_buf <= out23_bufn;
			out136_buf <= out136_bufn;
			out0_buf <= out0_bufn;
			out134_buf <= out134_bufn;
			out13_buf <= out13_bufn;
			out131_buf <= out131_bufn;
			out129_buf <= out129_bufn;
			out111_buf <= out111_bufn;
			out31_buf <= out31_bufn;
			out126_buf <= out126_bufn;
			out106_buf <= out106_bufn;
			out124_buf <= out124_bufn;
			out138_buf <= out138_bufn;
			out141_buf <= out141_bufn;
			out143_buf <= out143_bufn;
			out146_buf <= out146_bufn;
			out150_buf <= out150_bufn;
			out153_buf <= out153_bufn;
			out155_buf <= out155_bufn;
			out158_buf <= out158_bufn;
			out162_buf <= out162_bufn;
			out165_buf <= out165_bufn;
			out168_buf <= out168_bufn;
			out171_buf <= out171_bufn;
			out174_buf <= out174_bufn;
			out178_buf <= out178_bufn;
			out181_buf <= out181_bufn;
			out183_buf <= out183_bufn;
			out197_buf <= out197_bufn;
			out201_buf <= out201_bufn;
			out204_buf <= out204_bufn;
			out207_buf <= out207_bufn;
			out210_buf <= out210_bufn;
			out213_buf <= out213_bufn;
			out217_buf <= out217_bufn;
			out220_buf <= out220_bufn;
			out222_buf <= out222_bufn;
			out225_buf <= out225_bufn;
			out229_buf <= out229_bufn;
			out232_buf <= out232_bufn;
			out235_buf <= out235_bufn;
			out238_buf <= out238_bufn;
			out241_buf <= out241_bufn;
			out245_buf <= out245_bufn;
			out248_buf <= out248_bufn;
			out250_buf <= out250_bufn;
			out253_buf <= out253_bufn;
			out257_buf <= out257_bufn;
			out260_buf <= out260_bufn;
			out263_buf <= out263_bufn;
			out266_buf <= out266_bufn;
			out269_buf <= out269_bufn;
			out273_buf <= out273_bufn;
			out276_buf <= out276_bufn;
			out278_buf <= out278_bufn;
			out280_buf <= out280_bufn;
			out281_buf <= out281_bufn;
			out282_buf <= out282_bufn;
			out284_buf <= out284_bufn;
			out285_buf <= out285_bufn;
			out287_buf <= out287_bufn;
			out288_buf <= out288_bufn;
			out289_buf <= out289_bufn;
			out290_buf <= out290_bufn;
			out291_buf <= out291_bufn;
			out292_buf <= out292_bufn;
			out293_buf <= out293_bufn;
			out294_buf <= out294_bufn;
			out295_buf <= out295_bufn;
			out296_buf <= out296_bufn;
			out312_buf <= out312_bufn;
			out313_buf <= out313_bufn;
			out314_buf <= out314_bufn;
			out315_buf <= out315_bufn;
			out318_buf <= out318_bufn;
			out322_buf <= out322_bufn;
			out323_buf <= out323_bufn;
			out324_buf <= out324_bufn;
			out325_buf <= out325_bufn;
			out326_buf <= out326_bufn;
			out327_buf <= out327_bufn;
			out328_buf <= out328_bufn;
			out333_buf <= out333_bufn;
			out341_buf <= out341_bufn;
			out342_buf <= out342_bufn;
			out343_buf <= out343_bufn;
			out344_buf <= out344_bufn;
			out346_buf <= out346_bufn;
			out349_buf <= out349_bufn;
			out351_buf <= out351_bufn;
			out352_buf <= out352_bufn;
			out353_buf <= out353_bufn;
			out354_buf <= out354_bufn;
			out357_buf <= out357_bufn;
			out361_buf <= out361_bufn;
			out364_buf <= out364_bufn;
			out366_buf <= out366_bufn;
			out371_buf <= out371_bufn;
			out393_buf <= out393_bufn;
			out394_buf <= out394_bufn;
			out395_buf <= out395_bufn;
			out400_buf <= out400_bufn;
			out401_buf <= out401_bufn;
			out404_buf <= out404_bufn;
			out407_buf <= out407_bufn;
			out408_buf <= out408_bufn;
			out409_buf <= out409_bufn;
			out410_buf <= out410_bufn;
			out413_buf <= out413_bufn;
			out414_buf <= out414_bufn;
			out417_buf <= out417_bufn;
			out418_buf <= out418_bufn;
			out422_buf <= out422_bufn;
			out426_buf <= out426_bufn;
			out428_buf <= out428_bufn;
			out431_buf <= out431_bufn;
			out433_buf <= out433_bufn;
			out434_buf <= out434_bufn;
			out435_buf <= out435_bufn;
			out436_buf <= out436_bufn;
			out437_buf <= out437_bufn;
			out438_buf <= out438_bufn;
			out440_buf <= out440_bufn;
			out444_buf <= out444_bufn;
			out446_buf <= out446_bufn;
			out451_buf <= out451_bufn;
			out457_buf <= out457_bufn;
			out458_buf <= out458_bufn;
			out459_buf <= out459_bufn;
			out460_buf <= out460_bufn;
			out461_buf <= out461_bufn;
			out463_buf <= out463_bufn;
			out464_buf <= out464_bufn;
			out466_buf <= out466_bufn;
			out468_buf <= out468_bufn;
			out472_buf <= out472_bufn;
			out475_buf <= out475_bufn;
			out481_buf <= out481_bufn;
			out482_buf <= out482_bufn;
			out483_buf <= out483_bufn;
			out487_buf <= out487_bufn;
			out495_buf <= out495_bufn;
			out496_buf <= out496_bufn;
			out497_buf <= out497_bufn;
			out499_buf <= out499_bufn;
			out500_buf <= out500_bufn;
			out512_buf <= out512_bufn;
			out517_buf <= out517_bufn;
			out518_buf <= out518_bufn;
			out521_buf <= out521_bufn;
			out524_buf <= out524_bufn;
			out525_buf <= out525_bufn;
			out526_buf <= out526_bufn;
			out531_buf <= out531_bufn;
			out554_buf <= out554_bufn;
			out562_buf <= out562_bufn;
			out566_buf <= out566_bufn;
			-- Retiming: counters
			rtmcounter0 <= rtmcounter0_next;
			-- Function calls: return IDs

		end if;
	end process;

	-- Combinatorial process
	-- Compute the next state
	-- Compute the outputs

	process (
		-- Inputs of the FSM
		reset, in0, in2, in3, in4, in5, in1, in6, in11, in7, in8, in9, in10,
		-- Retiming: outputs of the comparators
		rtmcmp90, rtmcmp95, rtmcmp98, rtmcmp104, rtmcmp148, rtmcmp167, rtmcmp174, rtmcmp181, rtmcmp183, rtmcmp194, rtmcmp197, rtmcmp203, rtmcmp205, rtmcmp215,
		-- Retiming: the counters
		rtmcounter0,
		-- Function calls: return IDs
		-- Current state
		state_cur
	)
	begin

		-- Reset the next state value

		state_next <= (others => '0');

		-- Default value to the outputs or output buffers

		out22 <= '0';
		out4 <= '0';
		out122_bufn <= '0';
		out50 <= '0';
		out121 <= '0';
		out36_bufn <= '0';
		out49_bufn <= '0';
		out35_bufn <= '0';
		out99 <= '0';
		out52 <= '0';
		out18 <= '0';
		out33 <= '0';
		out123 <= '0';
		out101 <= '0';
		out90 <= '0';
		out91 <= '0';
		out27_bufn <= '0';
		out16_bufn <= '0';
		out26 <= '0';
		out21 <= '0';
		out24 <= '0';
		out54 <= '0';
		out25_bufn <= '0';
		out20_bufn <= '0';
		out58 <= '0';
		out30 <= '0';
		out8 <= '0';
		out57_bufn <= '0';
		out48 <= '0';
		out56 <= '0';
		out23_bufn <= '0';
		out29 <= '0';
		out19 <= '0';
		out136_bufn <= '0';
		out2 <= '0';
		out1 <= '0';
		out46 <= '0';
		out0_bufn <= '0';
		out135 <= '0';
		out118 <= '0';
		out116 <= '0';
		out14 <= '0';
		out134_bufn <= '0';
		out28 <= '0';
		out13_bufn <= '0';
		out133 <= '0';
		out131_bufn <= '0';
		out132 <= '0';
		out114 <= '0';
		out130 <= '0';
		out112 <= '0';
		out38 <= '0';
		out44 <= '0';
		out97 <= '0';
		out129_bufn <= '0';
		out111_bufn <= '0';
		out31_bufn <= '0';
		out126_bufn <= '0';
		out107 <= '0';
		out108 <= '0';
		out105 <= '0';
		out106_bufn <= '0';
		out125 <= '0';
		out120 <= '0';
		out124_bufn <= '0';
		out103 <= '0';
		out42 <= '0';
		out40 <= '0';
		out60 <= '0';
		out137 <= '0';
		out138_bufn <= '0';
		out140 <= '0';
		out141_bufn <= '0';
		out142 <= '0';
		out143_bufn <= '0';
		out145 <= '0';
		out146_bufn <= '0';
		out148 <= '0';
		out150_bufn <= '0';
		out153_bufn <= '0';
		out154 <= '0';
		out155_bufn <= '0';
		out156 <= '0';
		out157 <= '0';
		out158_bufn <= '0';
		out159 <= '0';
		out160 <= '0';
		out161 <= '0';
		out162_bufn <= '0';
		out164 <= '0';
		out165_bufn <= '0';
		out167 <= '0';
		out168_bufn <= '0';
		out170 <= '0';
		out171_bufn <= '0';
		out173 <= '0';
		out174_bufn <= '0';
		out176 <= '0';
		out178_bufn <= '0';
		out181_bufn <= '0';
		out182 <= '0';
		out183_bufn <= '0';
		out184 <= '0';
		out185 <= '0';
		out186 <= '0';
		out187 <= '0';
		out190 <= '0';
		out195 <= '0';
		out197_bufn <= '0';
		out198 <= '0';
		out199 <= '0';
		out200 <= '0';
		out201_bufn <= '0';
		out203 <= '0';
		out204_bufn <= '0';
		out206 <= '0';
		out207_bufn <= '0';
		out209 <= '0';
		out210_bufn <= '0';
		out212 <= '0';
		out213_bufn <= '0';
		out215 <= '0';
		out217_bufn <= '0';
		out220_bufn <= '0';
		out221 <= '0';
		out222_bufn <= '0';
		out223 <= '0';
		out224 <= '0';
		out225_bufn <= '0';
		out226 <= '0';
		out227 <= '0';
		out228 <= '0';
		out229_bufn <= '0';
		out231 <= '0';
		out232_bufn <= '0';
		out234 <= '0';
		out235_bufn <= '0';
		out237 <= '0';
		out238_bufn <= '0';
		out240 <= '0';
		out241_bufn <= '0';
		out243 <= '0';
		out245_bufn <= '0';
		out248_bufn <= '0';
		out249 <= '0';
		out250_bufn <= '0';
		out251 <= '0';
		out252 <= '0';
		out253_bufn <= '0';
		out254 <= '0';
		out255 <= '0';
		out256 <= '0';
		out257_bufn <= '0';
		out259 <= '0';
		out260_bufn <= '0';
		out262 <= '0';
		out263_bufn <= '0';
		out265 <= '0';
		out266_bufn <= '0';
		out268 <= '0';
		out269_bufn <= '0';
		out271 <= '0';
		out273_bufn <= '0';
		out276_bufn <= '0';
		out277 <= '0';
		out278_bufn <= '0';
		out279 <= '0';
		out280_bufn <= '0';
		out281_bufn <= '0';
		out282_bufn <= '0';
		out283 <= '0';
		out284_bufn <= '0';
		out285_bufn <= '0';
		out286 <= '0';
		out287_bufn <= '0';
		out288_bufn <= '0';
		out289_bufn <= '0';
		out290_bufn <= '0';
		out291_bufn <= '0';
		out292_bufn <= '0';
		out293_bufn <= '0';
		out294_bufn <= '0';
		out295_bufn <= '0';
		out296_bufn <= '0';
		out297 <= '0';
		out298 <= '0';
		out311 <= '0';
		out312_bufn <= '0';
		out313_bufn <= '0';
		out314_bufn <= '0';
		out315_bufn <= '0';
		out316 <= '0';
		out318_bufn <= '0';
		out321 <= '0';
		out322_bufn <= '0';
		out323_bufn <= '0';
		out324_bufn <= '0';
		out325_bufn <= '0';
		out326_bufn <= '0';
		out327_bufn <= '0';
		out328_bufn <= '0';
		out329 <= '0';
		out333_bufn <= '0';
		out341_bufn <= '0';
		out342_bufn <= '0';
		out343_bufn <= '0';
		out344_bufn <= '0';
		out345 <= '0';
		out346_bufn <= '0';
		out349_bufn <= '0';
		out350 <= '0';
		out351_bufn <= '0';
		out352_bufn <= '0';
		out353_bufn <= '0';
		out354_bufn <= '0';
		out355 <= '0';
		out357_bufn <= '0';
		out361_bufn <= '0';
		out362 <= '0';
		out363 <= '0';
		out364_bufn <= '0';
		out366_bufn <= '0';
		out367 <= '0';
		out371_bufn <= '0';
		out372 <= '0';
		out373 <= '0';
		out382 <= '0';
		out383 <= '0';
		out385 <= '0';
		out393_bufn <= '0';
		out394_bufn <= '0';
		out395_bufn <= '0';
		out396 <= '0';
		out398 <= '0';
		out400_bufn <= '0';
		out401_bufn <= '0';
		out402 <= '0';
		out404_bufn <= '0';
		out406 <= '0';
		out407_bufn <= '0';
		out408_bufn <= '0';
		out409_bufn <= '0';
		out410_bufn <= '0';
		out411 <= '0';
		out412 <= '0';
		out413_bufn <= '0';
		out414_bufn <= '0';
		out416 <= '0';
		out417_bufn <= '0';
		out418_bufn <= '0';
		out419 <= '0';
		out422_bufn <= '0';
		out423 <= '0';
		out425 <= '0';
		out426_bufn <= '0';
		out428_bufn <= '0';
		out429 <= '0';
		out430 <= '0';
		out431_bufn <= '0';
		out433_bufn <= '0';
		out434_bufn <= '0';
		out435_bufn <= '0';
		out436_bufn <= '0';
		out437_bufn <= '0';
		out438_bufn <= '0';
		out440_bufn <= '0';
		out441 <= '0';
		out443 <= '0';
		out444_bufn <= '0';
		out445 <= '0';
		out446_bufn <= '0';
		out447 <= '0';
		out450 <= '0';
		out451_bufn <= '0';
		out454 <= '0';
		out455 <= '0';
		out457_bufn <= '0';
		out458_bufn <= '0';
		out459_bufn <= '0';
		out460_bufn <= '0';
		out461_bufn <= '0';
		out462 <= '0';
		out463_bufn <= '0';
		out464_bufn <= '0';
		out465 <= '0';
		out466_bufn <= '0';
		out467 <= '0';
		out468_bufn <= '0';
		out469 <= '0';
		out472_bufn <= '0';
		out475_bufn <= '0';
		out481_bufn <= '0';
		out482_bufn <= '0';
		out483_bufn <= '0';
		out484 <= '0';
		out487_bufn <= '0';
		out488 <= '0';
		out491 <= '0';
		out495_bufn <= '0';
		out496_bufn <= '0';
		out497_bufn <= '0';
		out498 <= '0';
		out499_bufn <= '0';
		out500_bufn <= '0';
		out501 <= '0';
		out512_bufn <= '0';
		out513 <= '0';
		out517_bufn <= '0';
		out518_bufn <= '0';
		out519 <= '0';
		out521_bufn <= '0';
		out522 <= '0';
		out524_bufn <= '0';
		out525_bufn <= '0';
		out526_bufn <= '0';
		out527 <= '0';
		out528 <= '0';
		out531_bufn <= '0';
		out540 <= '0';
		out542 <= '0';
		out544 <= '0';
		out545 <= '0';
		out554_bufn <= '0';
		out555 <= '0';
		out559 <= '0';
		out560 <= '0';
		out561 <= '0';
		out562_bufn <= '0';
		out563 <= '0';
		out566_bufn <= '0';
		out567 <= '0';
		out570 <= '0';
		out572 <= '0';
		out575 <= '0';
		out577 <= '0';
		out578 <= '0';
		out580 <= '0';
		out581 <= '0';

		-- Retiming: default value for counters
		rtmcounter0_next <= (others => '0');

		-- Function calls: default values (no change)

		-- For all states, compute the next state bits
		--   And the outputs, and the next value for buffered outputs

		if state_cur(0) = '1' then
			-- Next state
			state_next(109) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out1 <= '1';
			out2 <= '1';
		end if;

		if state_cur(1) = '1' then
			-- Next state
			if (in0) = '1' then
				state_next(1) <= '1';
				-- Next values for buffered outputs
				out13_bufn <= '1';
			else
				-- Return from function: memextrct_0
				state_next(88) <= '1';
				-- Next values for buffered outputs
			end if;
			-- Assignment of non-buffered outputs
			out14 <= '1';
			out8 <= '1';
			out4 <= '1';
		end if;

		if state_cur(2) = '1' then
			-- Next state
			state_next(1) <= '1';
			-- Next values for buffered outputs
			out13_bufn <= '1';
			-- Assignment of non-buffered outputs
			out18 <= '1';
		end if;

		if state_cur(3) = '1' then
			-- Next state
			state_next(0) <= '1';
			-- Next values for buffered outputs
			out0_bufn <= '1';
			-- Assignment of non-buffered outputs
			out21 <= '1';
			out2 <= '1';
			out19 <= '1';
		end if;

		if state_cur(4) = '1' then
			-- Next state
			state_next(3) <= '1';
			-- Next values for buffered outputs
			out20_bufn <= '1';
			out0_bufn <= '1';
			-- Assignment of non-buffered outputs
			out21 <= '1';
			out2 <= '1';
			out22 <= '1';
		end if;

		if state_cur(5) = '1' then
			-- Next state
			state_next(4) <= '1';
			-- Next values for buffered outputs
			out23_bufn <= '1';
			out0_bufn <= '1';
			-- Assignment of non-buffered outputs
			out21 <= '1';
			out2 <= '1';
			out24 <= '1';
		end if;

		if state_cur(6) = '1' then
			-- Next state
			state_next(5) <= '1';
			-- Next values for buffered outputs
			out25_bufn <= '1';
			out0_bufn <= '1';
			-- Assignment of non-buffered outputs
			out21 <= '1';
			out2 <= '1';
			out26 <= '1';
		end if;

		-- Info: This is the init/reset state
		if state_cur(7) = '1' then
			-- Next state
			if (not (in2)) = '1' then
				state_next(7) <= '1';
				-- Next values for buffered outputs
			else
				if (in1) = '1' then
					state_next(60) <= '1';
					-- Next values for buffered outputs
				else
					state_next(154) <= '1';
					-- Next values for buffered outputs
				end if;
			end if;
			-- Assignment of non-buffered outputs
			out28 <= '1';
			out29 <= '1';
		end if;

		if state_cur(8) = '1' then
			-- Next state
			state_next(6) <= '1';
			-- Next values for buffered outputs
			out27_bufn <= '1';
			out0_bufn <= '1';
			-- Assignment of non-buffered outputs
			out21 <= '1';
			out2 <= '1';
			out30 <= '1';
		end if;

		if state_cur(9) = '1' then
			-- Next state
			state_next(9) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
		end if;

		if state_cur(10) = '1' then
			-- Next state
			state_next(8) <= '1';
			-- Next values for buffered outputs
			out31_bufn <= '1';
			out0_bufn <= '1';
			-- Assignment of non-buffered outputs
			out21 <= '1';
			out33 <= '1';
			out2 <= '1';
		end if;

		if state_cur(11) = '1' then
			-- Next state
			state_next(10) <= '1';
			-- Next values for buffered outputs
			out0_bufn <= '1';
			-- Assignment of non-buffered outputs
			out21 <= '1';
			out2 <= '1';
		end if;

		if state_cur(12) = '1' then
			-- Next state
			state_next(11) <= '1';
			-- Next values for buffered outputs
			out35_bufn <= '1';
			out0_bufn <= '1';
			-- Assignment of non-buffered outputs
			out21 <= '1';
		end if;

		if state_cur(13) = '1' then
			-- Next state
			state_next(12) <= '1';
			-- Next values for buffered outputs
			out36_bufn <= '1';
			-- Assignment of non-buffered outputs
			out52 <= '1';
			out50 <= '1';
			out48 <= '1';
			out46 <= '1';
			out44 <= '1';
			out42 <= '1';
			out40 <= '1';
			out38 <= '1';
		end if;

		if state_cur(14) = '1' then
			-- Next state
			state_next(13) <= '1';
			-- Next values for buffered outputs
			out49_bufn <= '1';
			-- Assignment of non-buffered outputs
			out60 <= '1';
			out58 <= '1';
			out56 <= '1';
			out54 <= '1';
		end if;

		if state_cur(15) = '1' then
			-- Next state
			if (in3) = '1' then
				state_next(15) <= '1';
				-- Next values for buffered outputs
				out13_bufn <= '1';
			else
				-- Return from function: memextrct_1
				state_next(88) <= '1';
				-- Next values for buffered outputs
			end if;
			-- Assignment of non-buffered outputs
			out14 <= '1';
			out91 <= '1';
			out90 <= '1';
		end if;

		if state_cur(16) = '1' then
			-- Next state
			if (in5) = '1' then
				-- Function call: memextrct_1
				state_next(19) <= '1';
				-- Next values for buffered outputs
				out16_bufn <= '1';
			else
				if (in4) = '1' then
					-- Function call: memextrct_0
					state_next(2) <= '1';
					-- Next values for buffered outputs
					out16_bufn <= '1';
				else
					state_next(88) <= '1';
					-- Next values for buffered outputs
				end if;
			end if;
			-- Assignment of non-buffered outputs
			out97 <= '1';
		end if;

		if state_cur(17) = '1' then
			-- Next state
			state_next(14) <= '1';
			-- Next values for buffered outputs
			out57_bufn <= '1';
			-- Assignment of non-buffered outputs
			out105 <= '1';
			out103 <= '1';
			out101 <= '1';
			out99 <= '1';
		end if;

		if state_cur(18) = '1' then
			-- Next state
			state_next(17) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out118 <= '1';
			out116 <= '1';
			out114 <= '1';
			out112 <= '1';
			out108 <= '1';
			out107 <= '1';
		end if;

		if state_cur(19) = '1' then
			-- Next state
			state_next(15) <= '1';
			-- Next values for buffered outputs
			out13_bufn <= '1';
			-- Assignment of non-buffered outputs
			out18 <= '1';
		end if;

		if state_cur(20) = '1' then
			-- Next state
			state_next(18) <= '1';
			-- Next values for buffered outputs
			out111_bufn <= '1';
			out106_bufn <= '1';
			-- Assignment of non-buffered outputs
			out52 <= '1';
			out21 <= '1';
			out125 <= '1';
			out123 <= '1';
			out108 <= '1';
			out121 <= '1';
		end if;

		if state_cur(21) = '1' then
			-- Next state
			state_next(20) <= '1';
			-- Next values for buffered outputs
			out126_bufn <= '1';
			out20_bufn <= '1';
			out124_bufn <= '1';
			out122_bufn <= '1';
			out106_bufn <= '1';
			-- Assignment of non-buffered outputs
			out132 <= '1';
			out50 <= '1';
			out21 <= '1';
			out130 <= '1';
			out108 <= '1';
		end if;

		if state_cur(22) = '1' then
			-- Next state
			state_next(21) <= '1';
			-- Next values for buffered outputs
			out131_bufn <= '1';
			out23_bufn <= '1';
			out129_bufn <= '1';
			out106_bufn <= '1';
			-- Assignment of non-buffered outputs
			out48 <= '1';
			out21 <= '1';
			out137 <= '1';
			out135 <= '1';
			out108 <= '1';
			out133 <= '1';
		end if;

		if state_cur(23) = '1' then
			-- Next state
			state_next(22) <= '1';
			-- Next values for buffered outputs
			out138_bufn <= '1';
			out25_bufn <= '1';
			out136_bufn <= '1';
			out134_bufn <= '1';
			out106_bufn <= '1';
			-- Assignment of non-buffered outputs
			out46 <= '1';
			out21 <= '1';
			out142 <= '1';
			out140 <= '1';
			out108 <= '1';
		end if;

		if state_cur(24) = '1' then
			-- Next state
			state_next(23) <= '1';
			-- Next values for buffered outputs
			out143_bufn <= '1';
			out27_bufn <= '1';
			out141_bufn <= '1';
			out106_bufn <= '1';
			-- Assignment of non-buffered outputs
			out44 <= '1';
			out21 <= '1';
			out145 <= '1';
			out108 <= '1';
		end if;

		if state_cur(25) = '1' then
			-- Next state
			state_next(24) <= '1';
			-- Next values for buffered outputs
			out146_bufn <= '1';
			out31_bufn <= '1';
			out106_bufn <= '1';
			-- Assignment of non-buffered outputs
			out42 <= '1';
			out21 <= '1';
			out148 <= '1';
			out108 <= '1';
		end if;

		if state_cur(26) = '1' then
			-- Next state
			state_next(25) <= '1';
			-- Next values for buffered outputs
			out150_bufn <= '1';
			out106_bufn <= '1';
			-- Assignment of non-buffered outputs
			out154 <= '1';
			out40 <= '1';
			out21 <= '1';
			out108 <= '1';
		end if;

		if state_cur(27) = '1' then
			-- Next state
			state_next(26) <= '1';
			-- Next values for buffered outputs
			out153_bufn <= '1';
			out35_bufn <= '1';
			out106_bufn <= '1';
			-- Assignment of non-buffered outputs
			out156 <= '1';
			out38 <= '1';
			out21 <= '1';
		end if;

		if state_cur(28) = '1' then
			-- Next state
			state_next(27) <= '1';
			-- Next values for buffered outputs
			out155_bufn <= '1';
			out36_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out46 <= '1';
			out52 <= '1';
			out48 <= '1';
			out44 <= '1';
			out42 <= '1';
			out40 <= '1';
			out38 <= '1';
		end if;

		if state_cur(29) = '1' then
			-- Next state
			state_next(28) <= '1';
			-- Next values for buffered outputs
			out49_bufn <= '1';
			-- Assignment of non-buffered outputs
			out60 <= '1';
			out157 <= '1';
			out58 <= '1';
			out56 <= '1';
			out54 <= '1';
		end if;

		if state_cur(30) = '1' then
			-- Next state
			state_next(29) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out105 <= '1';
			out103 <= '1';
			out101 <= '1';
			out99 <= '1';
		end if;

		if state_cur(31) = '1' then
			-- Next state
			state_next(30) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out118 <= '1';
			out116 <= '1';
			out114 <= '1';
			out112 <= '1';
			out160 <= '1';
			out159 <= '1';
		end if;

		if state_cur(32) = '1' then
			-- Next state
			state_next(31) <= '1';
			-- Next values for buffered outputs
			out111_bufn <= '1';
			out158_bufn <= '1';
			-- Assignment of non-buffered outputs
			out52 <= '1';
			out21 <= '1';
			out125 <= '1';
			out123 <= '1';
			out161 <= '1';
			out160 <= '1';
		end if;

		if state_cur(33) = '1' then
			-- Next state
			state_next(32) <= '1';
			-- Next values for buffered outputs
			out162_bufn <= '1';
			out20_bufn <= '1';
			out124_bufn <= '1';
			out122_bufn <= '1';
			out158_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out21 <= '1';
			out130 <= '1';
			out164 <= '1';
			out160 <= '1';
		end if;

		if state_cur(34) = '1' then
			-- Next state
			state_next(33) <= '1';
			-- Next values for buffered outputs
			out165_bufn <= '1';
			out23_bufn <= '1';
			out129_bufn <= '1';
			out158_bufn <= '1';
			-- Assignment of non-buffered outputs
			out48 <= '1';
			out21 <= '1';
			out137 <= '1';
			out135 <= '1';
			out167 <= '1';
			out160 <= '1';
		end if;

		if state_cur(35) = '1' then
			-- Next state
			state_next(34) <= '1';
			-- Next values for buffered outputs
			out168_bufn <= '1';
			out25_bufn <= '1';
			out136_bufn <= '1';
			out134_bufn <= '1';
			out158_bufn <= '1';
			-- Assignment of non-buffered outputs
			out46 <= '1';
			out21 <= '1';
			out142 <= '1';
			out170 <= '1';
			out160 <= '1';
		end if;

		if state_cur(36) = '1' then
			-- Next state
			state_next(35) <= '1';
			-- Next values for buffered outputs
			out171_bufn <= '1';
			out27_bufn <= '1';
			out141_bufn <= '1';
			out158_bufn <= '1';
			-- Assignment of non-buffered outputs
			out44 <= '1';
			out21 <= '1';
			out173 <= '1';
			out160 <= '1';
		end if;

		if state_cur(37) = '1' then
			-- Next state
			state_next(36) <= '1';
			-- Next values for buffered outputs
			out174_bufn <= '1';
			out31_bufn <= '1';
			out158_bufn <= '1';
			-- Assignment of non-buffered outputs
			out42 <= '1';
			out21 <= '1';
			out176 <= '1';
			out160 <= '1';
		end if;

		if state_cur(38) = '1' then
			-- Next state
			state_next(37) <= '1';
			-- Next values for buffered outputs
			out178_bufn <= '1';
			out158_bufn <= '1';
			-- Assignment of non-buffered outputs
			out182 <= '1';
			out40 <= '1';
			out21 <= '1';
			out160 <= '1';
		end if;

		if state_cur(39) = '1' then
			-- Next state
			state_next(38) <= '1';
			-- Next values for buffered outputs
			out181_bufn <= '1';
			out35_bufn <= '1';
			out158_bufn <= '1';
			-- Assignment of non-buffered outputs
			out184 <= '1';
			out38 <= '1';
			out21 <= '1';
		end if;

		if state_cur(40) = '1' then
			-- Next state
			state_next(39) <= '1';
			-- Next values for buffered outputs
			out183_bufn <= '1';
			out36_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out46 <= '1';
			out52 <= '1';
			out48 <= '1';
			out44 <= '1';
			out42 <= '1';
			out40 <= '1';
			out38 <= '1';
		end if;

		if state_cur(41) = '1' then
			-- Next state
			state_next(40) <= '1';
			-- Next values for buffered outputs
			out49_bufn <= '1';
			-- Assignment of non-buffered outputs
			out60 <= '1';
			out185 <= '1';
			out58 <= '1';
			out56 <= '1';
			out54 <= '1';
		end if;

		if state_cur(42) = '1' then
			-- Next state
			state_next(41) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out105 <= '1';
			out103 <= '1';
			out101 <= '1';
			out99 <= '1';
		end if;

		if state_cur(43) = '1' then
			-- Next state
			if (in7) = '1' then
				state_next(60) <= '1';
				-- Next values for buffered outputs
			else
				if (not (in6)) = '1' then
					state_next(43) <= '1';
					-- Next values for buffered outputs
				else
					state_next(108) <= '1';
					-- Next values for buffered outputs
					out371_bufn <= '1';
				end if;
			end if;
			-- Assignment of non-buffered outputs
			out190 <= '1';
			out187 <= '1';
			out186 <= '1';
		end if;

		if state_cur(44) = '1' then
			-- Next state
			if (in7) = '1' then
				state_next(60) <= '1';
				-- Next values for buffered outputs
			else
				if (not (in8)) = '1' then
					state_next(44) <= '1';
					-- Next values for buffered outputs
				else
					state_next(110) <= '1';
					-- Next values for buffered outputs
					out371_bufn <= '1';
				end if;
			end if;
			-- Assignment of non-buffered outputs
			out195 <= '1';
			out187 <= '1';
		end if;

		if state_cur(45) = '1' then
			-- Next state
			state_next(42) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out118 <= '1';
			out116 <= '1';
			out114 <= '1';
			out112 <= '1';
			out199 <= '1';
			out198 <= '1';
		end if;

		if state_cur(46) = '1' then
			-- Next state
			state_next(45) <= '1';
			-- Next values for buffered outputs
			out111_bufn <= '1';
			out197_bufn <= '1';
			-- Assignment of non-buffered outputs
			out52 <= '1';
			out21 <= '1';
			out125 <= '1';
			out123 <= '1';
			out200 <= '1';
			out199 <= '1';
		end if;

		if state_cur(47) = '1' then
			-- Next state
			state_next(46) <= '1';
			-- Next values for buffered outputs
			out201_bufn <= '1';
			out20_bufn <= '1';
			out124_bufn <= '1';
			out122_bufn <= '1';
			out197_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out21 <= '1';
			out130 <= '1';
			out203 <= '1';
			out199 <= '1';
		end if;

		if state_cur(48) = '1' then
			-- Next state
			state_next(47) <= '1';
			-- Next values for buffered outputs
			out204_bufn <= '1';
			out23_bufn <= '1';
			out129_bufn <= '1';
			out197_bufn <= '1';
			-- Assignment of non-buffered outputs
			out48 <= '1';
			out21 <= '1';
			out137 <= '1';
			out135 <= '1';
			out206 <= '1';
			out199 <= '1';
		end if;

		if state_cur(49) = '1' then
			-- Next state
			state_next(48) <= '1';
			-- Next values for buffered outputs
			out207_bufn <= '1';
			out25_bufn <= '1';
			out136_bufn <= '1';
			out134_bufn <= '1';
			out197_bufn <= '1';
			-- Assignment of non-buffered outputs
			out46 <= '1';
			out21 <= '1';
			out142 <= '1';
			out209 <= '1';
			out199 <= '1';
		end if;

		if state_cur(50) = '1' then
			-- Next state
			state_next(49) <= '1';
			-- Next values for buffered outputs
			out210_bufn <= '1';
			out27_bufn <= '1';
			out141_bufn <= '1';
			out197_bufn <= '1';
			-- Assignment of non-buffered outputs
			out44 <= '1';
			out21 <= '1';
			out212 <= '1';
			out199 <= '1';
		end if;

		if state_cur(51) = '1' then
			-- Next state
			state_next(50) <= '1';
			-- Next values for buffered outputs
			out213_bufn <= '1';
			out31_bufn <= '1';
			out197_bufn <= '1';
			-- Assignment of non-buffered outputs
			out42 <= '1';
			out21 <= '1';
			out215 <= '1';
			out199 <= '1';
		end if;

		if state_cur(52) = '1' then
			-- Next state
			state_next(51) <= '1';
			-- Next values for buffered outputs
			out217_bufn <= '1';
			out197_bufn <= '1';
			-- Assignment of non-buffered outputs
			out221 <= '1';
			out40 <= '1';
			out21 <= '1';
			out199 <= '1';
		end if;

		if state_cur(53) = '1' then
			-- Next state
			state_next(52) <= '1';
			-- Next values for buffered outputs
			out220_bufn <= '1';
			out35_bufn <= '1';
			out197_bufn <= '1';
			-- Assignment of non-buffered outputs
			out223 <= '1';
			out38 <= '1';
			out21 <= '1';
		end if;

		if state_cur(54) = '1' then
			-- Next state
			state_next(53) <= '1';
			-- Next values for buffered outputs
			out222_bufn <= '1';
			out36_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out46 <= '1';
			out52 <= '1';
			out48 <= '1';
			out44 <= '1';
			out42 <= '1';
			out40 <= '1';
			out38 <= '1';
		end if;

		if state_cur(55) = '1' then
			-- Next state
			state_next(54) <= '1';
			-- Next values for buffered outputs
			out49_bufn <= '1';
			-- Assignment of non-buffered outputs
			out60 <= '1';
			out224 <= '1';
			out58 <= '1';
			out56 <= '1';
			out54 <= '1';
		end if;

		if state_cur(56) = '1' then
			-- Next state
			state_next(55) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out105 <= '1';
			out103 <= '1';
			out101 <= '1';
			out99 <= '1';
		end if;

		if state_cur(57) = '1' then
			-- Next state
			state_next(56) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out118 <= '1';
			out116 <= '1';
			out114 <= '1';
			out112 <= '1';
			out227 <= '1';
			out226 <= '1';
		end if;

		if state_cur(58) = '1' then
			-- Next state
			state_next(57) <= '1';
			-- Next values for buffered outputs
			out111_bufn <= '1';
			out225_bufn <= '1';
			-- Assignment of non-buffered outputs
			out52 <= '1';
			out21 <= '1';
			out125 <= '1';
			out123 <= '1';
			out228 <= '1';
			out227 <= '1';
		end if;

		if state_cur(59) = '1' then
			-- Next state
			state_next(58) <= '1';
			-- Next values for buffered outputs
			out229_bufn <= '1';
			out20_bufn <= '1';
			out124_bufn <= '1';
			out122_bufn <= '1';
			out225_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out21 <= '1';
			out130 <= '1';
			out231 <= '1';
			out227 <= '1';
		end if;

		if state_cur(60) = '1' then
			-- Next state
			state_next(87) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out18 <= '1';
		end if;

		if state_cur(61) = '1' then
			-- Next state
			state_next(59) <= '1';
			-- Next values for buffered outputs
			out232_bufn <= '1';
			out23_bufn <= '1';
			out129_bufn <= '1';
			out225_bufn <= '1';
			-- Assignment of non-buffered outputs
			out48 <= '1';
			out21 <= '1';
			out137 <= '1';
			out135 <= '1';
			out234 <= '1';
			out227 <= '1';
		end if;

		if state_cur(62) = '1' then
			-- Next state
			state_next(61) <= '1';
			-- Next values for buffered outputs
			out235_bufn <= '1';
			out25_bufn <= '1';
			out136_bufn <= '1';
			out134_bufn <= '1';
			out225_bufn <= '1';
			-- Assignment of non-buffered outputs
			out46 <= '1';
			out21 <= '1';
			out142 <= '1';
			out237 <= '1';
			out227 <= '1';
		end if;

		if state_cur(63) = '1' then
			-- Next state
			state_next(62) <= '1';
			-- Next values for buffered outputs
			out238_bufn <= '1';
			out27_bufn <= '1';
			out141_bufn <= '1';
			out225_bufn <= '1';
			-- Assignment of non-buffered outputs
			out44 <= '1';
			out21 <= '1';
			out240 <= '1';
			out227 <= '1';
		end if;

		if state_cur(64) = '1' then
			-- Next state
			state_next(63) <= '1';
			-- Next values for buffered outputs
			out241_bufn <= '1';
			out31_bufn <= '1';
			out225_bufn <= '1';
			-- Assignment of non-buffered outputs
			out42 <= '1';
			out21 <= '1';
			out243 <= '1';
			out227 <= '1';
		end if;

		if state_cur(65) = '1' then
			-- Next state
			state_next(64) <= '1';
			-- Next values for buffered outputs
			out245_bufn <= '1';
			out225_bufn <= '1';
			-- Assignment of non-buffered outputs
			out249 <= '1';
			out40 <= '1';
			out21 <= '1';
			out227 <= '1';
		end if;

		if state_cur(66) = '1' then
			-- Next state
			state_next(65) <= '1';
			-- Next values for buffered outputs
			out248_bufn <= '1';
			out35_bufn <= '1';
			out225_bufn <= '1';
			-- Assignment of non-buffered outputs
			out251 <= '1';
			out38 <= '1';
			out21 <= '1';
		end if;

		if state_cur(67) = '1' then
			-- Next state
			state_next(66) <= '1';
			-- Next values for buffered outputs
			out250_bufn <= '1';
			out36_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out46 <= '1';
			out52 <= '1';
			out48 <= '1';
			out44 <= '1';
			out42 <= '1';
			out40 <= '1';
			out38 <= '1';
		end if;

		if state_cur(68) = '1' then
			-- Next state
			state_next(67) <= '1';
			-- Next values for buffered outputs
			out49_bufn <= '1';
			-- Assignment of non-buffered outputs
			out60 <= '1';
			out252 <= '1';
			out58 <= '1';
			out56 <= '1';
			out54 <= '1';
		end if;

		if state_cur(69) = '1' then
			-- Next state
			state_next(68) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out105 <= '1';
			out103 <= '1';
			out101 <= '1';
			out99 <= '1';
		end if;

		if state_cur(70) = '1' then
			-- Next state
			state_next(69) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out118 <= '1';
			out116 <= '1';
			out114 <= '1';
			out112 <= '1';
			out255 <= '1';
			out254 <= '1';
		end if;

		if state_cur(71) = '1' then
			-- Next state
			state_next(70) <= '1';
			-- Next values for buffered outputs
			out111_bufn <= '1';
			out253_bufn <= '1';
			-- Assignment of non-buffered outputs
			out52 <= '1';
			out21 <= '1';
			out125 <= '1';
			out123 <= '1';
			out256 <= '1';
			out255 <= '1';
		end if;

		if state_cur(72) = '1' then
			-- Next state
			state_next(71) <= '1';
			-- Next values for buffered outputs
			out257_bufn <= '1';
			out20_bufn <= '1';
			out124_bufn <= '1';
			out122_bufn <= '1';
			out253_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out21 <= '1';
			out130 <= '1';
			out259 <= '1';
			out255 <= '1';
		end if;

		if state_cur(73) = '1' then
			-- Next state
			state_next(72) <= '1';
			-- Next values for buffered outputs
			out260_bufn <= '1';
			out23_bufn <= '1';
			out129_bufn <= '1';
			out253_bufn <= '1';
			-- Assignment of non-buffered outputs
			out48 <= '1';
			out21 <= '1';
			out137 <= '1';
			out135 <= '1';
			out262 <= '1';
			out255 <= '1';
		end if;

		if state_cur(74) = '1' then
			-- Next state
			state_next(73) <= '1';
			-- Next values for buffered outputs
			out263_bufn <= '1';
			out25_bufn <= '1';
			out136_bufn <= '1';
			out134_bufn <= '1';
			out253_bufn <= '1';
			-- Assignment of non-buffered outputs
			out46 <= '1';
			out21 <= '1';
			out142 <= '1';
			out265 <= '1';
			out255 <= '1';
		end if;

		if state_cur(75) = '1' then
			-- Next state
			state_next(74) <= '1';
			-- Next values for buffered outputs
			out266_bufn <= '1';
			out27_bufn <= '1';
			out141_bufn <= '1';
			out253_bufn <= '1';
			-- Assignment of non-buffered outputs
			out44 <= '1';
			out21 <= '1';
			out268 <= '1';
			out255 <= '1';
		end if;

		if state_cur(76) = '1' then
			-- Next state
			state_next(75) <= '1';
			-- Next values for buffered outputs
			out269_bufn <= '1';
			out31_bufn <= '1';
			out253_bufn <= '1';
			-- Assignment of non-buffered outputs
			out42 <= '1';
			out21 <= '1';
			out271 <= '1';
			out255 <= '1';
		end if;

		if state_cur(77) = '1' then
			-- Next state
			state_next(76) <= '1';
			-- Next values for buffered outputs
			out273_bufn <= '1';
			out253_bufn <= '1';
			-- Assignment of non-buffered outputs
			out277 <= '1';
			out40 <= '1';
			out21 <= '1';
			out255 <= '1';
		end if;

		if state_cur(78) = '1' then
			-- Next state
			state_next(77) <= '1';
			-- Next values for buffered outputs
			out276_bufn <= '1';
			out35_bufn <= '1';
			out253_bufn <= '1';
			-- Assignment of non-buffered outputs
			out279 <= '1';
			out38 <= '1';
			out21 <= '1';
		end if;

		if state_cur(79) = '1' then
			-- Next state
			state_next(80) <= '1';
			-- Next values for buffered outputs
			out285_bufn <= '1';
			out284_bufn <= '1';
			out269_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(80) = '1' then
			-- Next state
			state_next(113) <= '1';
			-- Next values for buffered outputs
			out395_bufn <= '1';
			out284_bufn <= '1';
			out146_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(81) = '1' then
			-- Next state
			state_next(82) <= '1';
			-- Next values for buffered outputs
			out290_bufn <= '1';
			out289_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(82) = '1' then
			-- Next state
			state_next(83) <= '1';
			-- Next values for buffered outputs
			out57_bufn <= '1';
			out292_bufn <= '1';
			out291_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(83) = '1' then
			-- Next state
			state_next(85) <= '1';
			-- Next values for buffered outputs
			out295_bufn <= '1';
			out294_bufn <= '1';
			-- Assignment of non-buffered outputs
			out58 <= '1';
			out118 <= '1';
			out286 <= '1';
		end if;

		if state_cur(84) = '1' then
			-- Next state
			state_next(89) <= '1';
			-- Next values for buffered outputs
			out313_bufn <= '1';
			out281_bufn <= '1';
			out312_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(85) = '1' then
			-- Next state
			state_next(86) <= '1';
			-- Next values for buffered outputs
			out296_bufn <= '1';
			out291_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(86) = '1' then
			-- Next state
			state_next(90) <= '1';
			-- Next values for buffered outputs
			out318_bufn <= '1';
			out280_bufn <= '1';
			out315_bufn <= '1';
			out314_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(87) = '1' then
			-- Next state
			if (in9) = '1' then
				state_next(87) <= '1';
				-- Next values for buffered outputs
			else
				state_next(16) <= '1';
				-- Next values for buffered outputs
				out16_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs
			out14 <= '1';
			out298 <= '1';
			out297 <= '1';
		end if;

		if state_cur(88) = '1' then
			-- Next state
			if (in1) = '1' then
				if (in5) = '1' then
					state_next(43) <= '1';
					-- Next values for buffered outputs
				else
					state_next(44) <= '1';
					-- Next values for buffered outputs
				end if;
			else
				state_next(9) <= '1';
				-- Next values for buffered outputs
			end if;
			-- Assignment of non-buffered outputs
			out311 <= '1';
		end if;

		if state_cur(89) = '1' then
			-- Next state
			state_next(112) <= '1';
			-- Next values for buffered outputs
			out394_bufn <= '1';
			out284_bufn <= '1';
			out393_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(90) = '1' then
			if rtmcmp90 = '1' then
				-- Next state
				state_next(93) <= '1';
				-- Next values for buffered outputs
				out57_bufn <= '1';
				out325_bufn <= '1';
				out324_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out103 <= '1';
				out105 <= '1';
				out56 <= '1';
				out137 <= '1';
				out125 <= '1';
				out116 <= '1';
				out283 <= '1';
			else  -- Stay in the current state
				state_next(90) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out318_bufn <= '1';
				out280_bufn <= '1';
				out315_bufn <= '1';
				out314_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out316 <= '1';
		end if;

		if state_cur(91) = '1' then
			-- Next state
			state_next(170) <= '1';
			-- Next values for buffered outputs
			out487_bufn <= '1';
			out284_bufn <= '1';
			out266_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
			out321 <= '1';
		end if;

		if state_cur(92) = '1' then
			-- Next state
			state_next(240) <= '1';
			-- Next values for buffered outputs
			out217_bufn <= '1';
			out295_bufn <= '1';
			out281_bufn <= '1';
			out562_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(93) = '1' then
			-- Next state
			state_next(101) <= '1';
			-- Next values for buffered outputs
			out323_bufn <= '1';
			out291_bufn <= '1';
			-- Assignment of non-buffered outputs
			out118 <= '1';
			out58 <= '1';
			out286 <= '1';
		end if;

		if state_cur(94) = '1' then
			-- Next state
			state_next(96) <= '1';
			-- Next values for buffered outputs
			out341_bufn <= '1';
			out281_bufn <= '1';
			out241_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(95) = '1' then
			if rtmcmp95 = '1' then
				-- Next state
				state_next(210) <= '1';
				-- Next values for buffered outputs
				out418_bufn <= '1';
				out351_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out130 <= '1';
				out101 <= '1';
				out142 <= '1';
				out112 <= '1';
				out99 <= '1';
				out54 <= '1';
				out123 <= '1';
				out135 <= '1';
				out114 <= '1';
				out286 <= '1';
			else  -- Stay in the current state
				state_next(95) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out333_bufn <= '1';
				out245_bufn <= '1';
				out318_bufn <= '1';
				out328_bufn <= '1';
				out327_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out329 <= '1';
		end if;

		if state_cur(96) = '1' then
			-- Next state
			state_next(91) <= '1';
			-- Next values for buffered outputs
			out322_bufn <= '1';
			out281_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(97) = '1' then
			-- Next state
			state_next(95) <= '1';
			-- Next values for buffered outputs
			out333_bufn <= '1';
			out245_bufn <= '1';
			out318_bufn <= '1';
			out328_bufn <= '1';
			out327_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(98) = '1' then
			if rtmcmp98 = '1' then
				-- Next state
				state_next(97) <= '1';
				-- Next values for buffered outputs
				out342_bufn <= '1';
				out324_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out125 <= '1';
				out137 <= '1';
				out116 <= '1';
				out56 <= '1';
				out283 <= '1';
			else  -- Stay in the current state
				state_next(98) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out346_bufn <= '1';
				out344_bufn <= '1';
				out312_bufn <= '1';
				out343_bufn <= '1';
				out314_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out345 <= '1';
		end if;

		if state_cur(99) = '1' then
			-- Next state
			state_next(119) <= '1';
			-- Next values for buffered outputs
			out36_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out46 <= '1';
			out52 <= '1';
			out48 <= '1';
			out44 <= '1';
			out42 <= '1';
			out40 <= '1';
			out38 <= '1';
		end if;

		if state_cur(100) = '1' then
			-- Next state
			state_next(233) <= '1';
			-- Next values for buffered outputs
			out566_bufn <= '1';
			out289_bufn <= '1';
			-- Assignment of non-buffered outputs
			out125 <= '1';
			out286 <= '1';
		end if;

		if state_cur(101) = '1' then
			-- Next state
			state_next(98) <= '1';
			-- Next values for buffered outputs
			out346_bufn <= '1';
			out344_bufn <= '1';
			out312_bufn <= '1';
			out343_bufn <= '1';
			out314_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(102) = '1' then
			-- Next state
			state_next(239) <= '1';
			-- Next values for buffered outputs
			out49_bufn <= '1';
			-- Assignment of non-buffered outputs
			out60 <= '1';
			out350 <= '1';
			out58 <= '1';
			out56 <= '1';
			out54 <= '1';
		end if;

		if state_cur(103) = '1' then
			-- Next state
			state_next(146) <= '1';
			-- Next values for buffered outputs
			out401_bufn <= '1';
			out444_bufn <= '1';
			out294_bufn <= '1';
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out60 <= '1';
			out283 <= '1';
		end if;

		if state_cur(104) = '1' then
			if rtmcmp104 = '1' then
				-- Next state
				state_next(103) <= '1';
				-- Next values for buffered outputs
				out352_bufn <= '1';
				out351_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out142 <= '1';
				out99 <= '1';
				out130 <= '1';
				out101 <= '1';
				out54 <= '1';
				out135 <= '1';
				out123 <= '1';
				out114 <= '1';
				out286 <= '1';
			else  -- Stay in the current state
				state_next(104) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out129_bufn <= '1';
				out357_bufn <= '1';
				out354_bufn <= '1';
				out353_bufn <= '1';
				out327_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out355 <= '1';
		end if;

		if state_cur(105) = '1' then
			-- Next state
			state_next(133) <= '1';
			-- Next values for buffered outputs
			out431_bufn <= '1';
			out23_bufn <= '1';
			out129_bufn <= '1';
			out361_bufn <= '1';
			-- Assignment of non-buffered outputs
			out48 <= '1';
			out21 <= '1';
			out137 <= '1';
			out135 <= '1';
			out363 <= '1';
			out362 <= '1';
		end if;

		if state_cur(106) = '1' then
			-- Next state
			state_next(186) <= '1';
			-- Next values for buffered outputs
			out518_bufn <= '1';
			out284_bufn <= '1';
			out153_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(107) = '1' then
			-- Next state
			state_next(148) <= '1';
			-- Next values for buffered outputs
			out446_bufn <= '1';
			out413_bufn <= '1';
			out281_bufn <= '1';
			out250_bufn <= '1';
			-- Assignment of non-buffered outputs
			out112 <= '1';
			out367 <= '1';
			out283 <= '1';
		end if;

		if state_cur(108) = '1' then
			-- Next state
			if (in10) = '1' then
				state_next(109) <= '1';
				-- Next values for buffered outputs
			else
				state_next(154) <= '1';
				-- Next values for buffered outputs
			end if;
			-- Assignment of non-buffered outputs
			out372 <= '1';
		end if;

		if state_cur(109) = '1' then
			-- Next state
			state_next(43) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out382 <= '1';
			out373 <= '1';
		end if;

		if state_cur(110) = '1' then
			-- Next state
			if (in11) = '1' then
				state_next(44) <= '1';
				-- Next values for buffered outputs
			else
				state_next(111) <= '1';
				-- Next values for buffered outputs
				out284_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs
			out372 <= '1';
			out385 <= '1';
			out383 <= '1';
		end if;

		if state_cur(111) = '1' then
			-- Next state
			state_next(153) <= '1';
			-- Next values for buffered outputs
			out422_bufn <= '1';
			out284_bufn <= '1';
			out278_bufn <= '1';
			-- Assignment of non-buffered outputs
			out372 <= '1';
			out286 <= '1';
		end if;

		if state_cur(112) = '1' then
			-- Next state
			state_next(94) <= '1';
			-- Next values for buffered outputs
			out326_bufn <= '1';
			out284_bufn <= '1';
			out210_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(113) = '1' then
			-- Next state
			state_next(160) <= '1';
			-- Next values for buffered outputs
			out461_bufn <= '1';
			out281_bufn <= '1';
			out178_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(114) = '1' then
			-- Next state
			state_next(196) <= '1';
			-- Next values for buffered outputs
			out328_bufn <= '1';
			out284_bufn <= '1';
			out155_bufn <= '1';
			-- Assignment of non-buffered outputs
			out142 <= '1';
			out396 <= '1';
			out286 <= '1';
		end if;

		if state_cur(115) = '1' then
			-- Next state
			state_next(105) <= '1';
			-- Next values for buffered outputs
			out364_bufn <= '1';
			out25_bufn <= '1';
			out136_bufn <= '1';
			out134_bufn <= '1';
			out361_bufn <= '1';
			-- Assignment of non-buffered outputs
			out46 <= '1';
			out21 <= '1';
			out142 <= '1';
			out398 <= '1';
			out363 <= '1';
		end if;

		if state_cur(116) = '1' then
			-- Next state
			state_next(120) <= '1';
			-- Next values for buffered outputs
			out407_bufn <= '1';
			out281_bufn <= '1';
			out168_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(117) = '1' then
			-- Next state
			state_next(211) <= '1';
			-- Next values for buffered outputs
			out458_bufn <= '1';
			out475_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(118) = '1' then
			-- Next state
			state_next(151) <= '1';
			-- Next values for buffered outputs
			out333_bufn <= '1';
			out31_bufn <= '1';
			out361_bufn <= '1';
			-- Assignment of non-buffered outputs
			out42 <= '1';
			out21 <= '1';
			out402 <= '1';
			out363 <= '1';
		end if;

		if state_cur(119) = '1' then
			-- Next state
			state_next(150) <= '1';
			-- Next values for buffered outputs
			out366_bufn <= '1';
			out35_bufn <= '1';
			out361_bufn <= '1';
			-- Assignment of non-buffered outputs
			out406 <= '1';
			out38 <= '1';
			out21 <= '1';
		end if;

		if state_cur(120) = '1' then
			-- Next state
			state_next(121) <= '1';
			-- Next values for buffered outputs
			out409_bufn <= '1';
			out281_bufn <= '1';
			out408_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(121) = '1' then
			-- Next state
			state_next(139) <= '1';
			-- Next values for buffered outputs
			out438_bufn <= '1';
			out284_bufn <= '1';
			out431_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(122) = '1' then
			-- Next state
			state_next(123) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out118 <= '1';
			out116 <= '1';
			out114 <= '1';
			out112 <= '1';
			out412 <= '1';
			out411 <= '1';
		end if;

		if state_cur(123) = '1' then
			-- Next state
			state_next(212) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out103 <= '1';
			out105 <= '1';
			out99 <= '1';
			out101 <= '1';
		end if;

		if state_cur(124) = '1' then
			-- Next state
			state_next(81) <= '1';
			-- Next values for buffered outputs
			out288_bufn <= '1';
			out287_bufn <= '1';
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out60 <= '1';
			out283 <= '1';
		end if;

		if state_cur(125) = '1' then
			-- Next state
			state_next(128) <= '1';
			-- Next values for buffered outputs
			out422_bufn <= '1';
			out287_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(126) = '1' then
			-- Next state
			state_next(125) <= '1';
			-- Next values for buffered outputs
			out414_bufn <= '1';
			out294_bufn <= '1';
			-- Assignment of non-buffered outputs
			out416 <= '1';
			out38 <= '1';
			out286 <= '1';
		end if;

		if state_cur(127) = '1' then
			-- Next state
			state_next(169) <= '1';
			-- Next values for buffered outputs
			out417_bufn <= '1';
			out483_bufn <= '1';
			out482_bufn <= '1';
			out318_bufn <= '1';
			-- Assignment of non-buffered outputs
			out112 <= '1';
			out419 <= '1';
			out283 <= '1';
		end if;

		if state_cur(128) = '1' then
			-- Next state
			state_next(124) <= '1';
			-- Next values for buffered outputs
			out413_bufn <= '1';
			out289_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(129) = '1' then
			-- Next state
			state_next(130) <= '1';
			-- Next values for buffered outputs
			out426_bufn <= '1';
			out27_bufn <= '1';
			out141_bufn <= '1';
			out410_bufn <= '1';
			-- Assignment of non-buffered outputs
			out44 <= '1';
			out21 <= '1';
			out423 <= '1';
			out412 <= '1';
		end if;

		if state_cur(130) = '1' then
			-- Next state
			state_next(143) <= '1';
			-- Next values for buffered outputs
			out435_bufn <= '1';
			out25_bufn <= '1';
			out136_bufn <= '1';
			out134_bufn <= '1';
			out410_bufn <= '1';
			-- Assignment of non-buffered outputs
			out46 <= '1';
			out21 <= '1';
			out142 <= '1';
			out425 <= '1';
			out412 <= '1';
		end if;

		if state_cur(131) = '1' then
			-- Next state
			state_next(102) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out103 <= '1';
			out105 <= '1';
			out99 <= '1';
			out101 <= '1';
		end if;

		if state_cur(132) = '1' then
			-- Next state
			state_next(144) <= '1';
			-- Next values for buffered outputs
			out111_bufn <= '1';
			-- Assignment of non-buffered outputs
			out114 <= '1';
			out429 <= '1';
			out52 <= '1';
			out286 <= '1';
		end if;

		if state_cur(133) = '1' then
			-- Next state
			state_next(237) <= '1';
			-- Next values for buffered outputs
			out475_bufn <= '1';
			out20_bufn <= '1';
			out124_bufn <= '1';
			out122_bufn <= '1';
			out361_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out21 <= '1';
			out130 <= '1';
			out430 <= '1';
			out363 <= '1';
		end if;

		if state_cur(134) = '1' then
			-- Next state
			state_next(227) <= '1';
			-- Next values for buffered outputs
			out496_bufn <= '1';
			out284_bufn <= '1';
			out263_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(135) = '1' then
			-- Next state
			state_next(117) <= '1';
			-- Next values for buffered outputs
			out352_bufn <= '1';
			out281_bufn <= '1';
			out401_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(136) = '1' then
			-- Next state
			state_next(135) <= '1';
			-- Next values for buffered outputs
			out434_bufn <= '1';
			out281_bufn <= '1';
			out165_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(137) = '1' then
			-- Next state
			state_next(228) <= '1';
			-- Next values for buffered outputs
			out463_bufn <= '1';
			out284_bufn <= '1';
			out260_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(138) = '1' then
			-- Next state
			state_next(137) <= '1';
			-- Next values for buffered outputs
			out436_bufn <= '1';
			out281_bufn <= '1';
			out435_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(139) = '1' then
			-- Next state
			state_next(229) <= '1';
			-- Next values for buffered outputs
			out495_bufn <= '1';
			out284_bufn <= '1';
			out204_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(140) = '1' then
			-- Next state
			state_next(126) <= '1';
			-- Next values for buffered outputs
			out324_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(141) = '1' then
			-- Next state
			state_next(142) <= '1';
			-- Next values for buffered outputs
			out122_bufn <= '1';
			out134_bufn <= '1';
			out400_bufn <= '1';
			out327_bufn <= '1';
			-- Assignment of non-buffered outputs
			out116 <= '1';
			out283 <= '1';
		end if;

		if state_cur(142) = '1' then
			-- Next state
			state_next(168) <= '1';
			-- Next values for buffered outputs
			out481_bufn <= '1';
			out351_bufn <= '1';
			-- Assignment of non-buffered outputs
			out54 <= '1';
			out123 <= '1';
			out135 <= '1';
			out114 <= '1';
			out286 <= '1';
		end if;

		if state_cur(143) = '1' then
			-- Next state
			state_next(149) <= '1';
			-- Next values for buffered outputs
			out451_bufn <= '1';
			out23_bufn <= '1';
			out129_bufn <= '1';
			out410_bufn <= '1';
			-- Assignment of non-buffered outputs
			out48 <= '1';
			out21 <= '1';
			out137 <= '1';
			out135 <= '1';
			out441 <= '1';
			out412 <= '1';
		end if;

		if state_cur(144) = '1' then
			-- Next state
			state_next(178) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out112 <= '1';
		end if;

		if state_cur(145) = '1' then
			-- Next state
			state_next(99) <= '1';
			-- Next values for buffered outputs
			out49_bufn <= '1';
			-- Assignment of non-buffered outputs
			out60 <= '1';
			out443 <= '1';
			out58 <= '1';
			out56 <= '1';
			out54 <= '1';
		end if;

		if state_cur(146) = '1' then
			-- Next state
			state_next(100) <= '1';
			-- Next values for buffered outputs
			out124_bufn <= '1';
			out349_bufn <= '1';
			out287_bufn <= '1';
			-- Assignment of non-buffered outputs
			out445 <= '1';
			out50 <= '1';
			out283 <= '1';
		end if;

		if state_cur(147) = '1' then
			-- Next state
			state_next(78) <= '1';
			-- Next values for buffered outputs
			out278_bufn <= '1';
			out36_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out46 <= '1';
			out52 <= '1';
			out48 <= '1';
			out44 <= '1';
			out42 <= '1';
			out40 <= '1';
			out38 <= '1';
		end if;

		if state_cur(148) = '1' then
			if rtmcmp148 = '1' then
				-- Next state
				state_next(172) <= '1';
				-- Next values for buffered outputs
				out296_bufn <= '1';
				out284_bufn <= '1';
				out220_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out103 <= '1';
				out125 <= '1';
				out99 <= '1';
				out123 <= '1';
				out283 <= '1';
			else  -- Stay in the current state
				state_next(148) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out446_bufn <= '1';
				out413_bufn <= '1';
				out281_bufn <= '1';
				out250_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out447 <= '1';
		end if;

		if state_cur(149) = '1' then
			-- Next state
			state_next(226) <= '1';
			-- Next values for buffered outputs
			out354_bufn <= '1';
			out20_bufn <= '1';
			out124_bufn <= '1';
			out122_bufn <= '1';
			out410_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out21 <= '1';
			out130 <= '1';
			out450 <= '1';
			out412 <= '1';
		end if;

		if state_cur(150) = '1' then
			-- Next state
			state_next(118) <= '1';
			-- Next values for buffered outputs
			out404_bufn <= '1';
			out361_bufn <= '1';
			-- Assignment of non-buffered outputs
			out454 <= '1';
			out40 <= '1';
			out21 <= '1';
			out363 <= '1';
		end if;

		if state_cur(151) = '1' then
			-- Next state
			state_next(115) <= '1';
			-- Next values for buffered outputs
			out393_bufn <= '1';
			out27_bufn <= '1';
			out141_bufn <= '1';
			out361_bufn <= '1';
			-- Assignment of non-buffered outputs
			out44 <= '1';
			out21 <= '1';
			out455 <= '1';
			out363 <= '1';
		end if;

		if state_cur(152) = '1' then
			-- Next state
			state_next(230) <= '1';
			-- Next values for buffered outputs
			out512_bufn <= '1';
			out281_bufn <= '1';
			out171_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(153) = '1' then
			-- Next state
			state_next(114) <= '1';
			-- Next values for buffered outputs
			out292_bufn <= '1';
			out284_bufn <= '1';
			out222_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(154) = '1' then
			-- Next state
			state_next(44) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out372 <= '1';
		end if;

		if state_cur(155) = '1' then
			-- Next state
			state_next(232) <= '1';
			-- Next values for buffered outputs
			out517_bufn <= '1';
			out284_bufn <= '1';
			out207_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(156) = '1' then
			-- Next state
			state_next(104) <= '1';
			-- Next values for buffered outputs
			out129_bufn <= '1';
			out357_bufn <= '1';
			out354_bufn <= '1';
			out353_bufn <= '1';
			out327_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(157) = '1' then
			-- Next state
			state_next(156) <= '1';
			-- Next values for buffered outputs
			out458_bufn <= '1';
			out324_bufn <= '1';
			-- Assignment of non-buffered outputs
			out56 <= '1';
			out137 <= '1';
			out116 <= '1';
			out283 <= '1';
		end if;

		if state_cur(158) = '1' then
			-- Next state
			state_next(157) <= '1';
			-- Next values for buffered outputs
			out136_bufn <= '1';
			out434_bufn <= '1';
			out314_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(159) = '1' then
			-- Next state
			state_next(158) <= '1';
			-- Next values for buffered outputs
			out459_bufn <= '1';
			out291_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(160) = '1' then
			-- Next state
			state_next(189) <= '1';
			-- Next values for buffered outputs
			out525_bufn <= '1';
			out281_bufn <= '1';
			out245_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(161) = '1' then
			-- Next state
			state_next(106) <= '1';
			-- Next values for buffered outputs
			out288_bufn <= '1';
			out284_bufn <= '1';
			out276_bufn <= '1';
			-- Assignment of non-buffered outputs
			out60 <= '1';
			out58 <= '1';
			out56 <= '1';
			out54 <= '1';
			out462 <= '1';
			out283 <= '1';
		end if;

		if state_cur(162) = '1' then
			-- Next state
			state_next(159) <= '1';
			-- Next values for buffered outputs
			out460_bufn <= '1';
			out289_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(163) = '1' then
			-- Next state
			state_next(162) <= '1';
			-- Next values for buffered outputs
			out463_bufn <= '1';
			out287_bufn <= '1';
			-- Assignment of non-buffered outputs
			out118 <= '1';
			out58 <= '1';
			out465 <= '1';
			out48 <= '1';
			out283 <= '1';
		end if;

		if state_cur(164) = '1' then
			-- Next state
			state_next(163) <= '1';
			-- Next values for buffered outputs
			out57_bufn <= '1';
			out408_bufn <= '1';
			out464_bufn <= '1';
			out294_bufn <= '1';
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out60 <= '1';
			out103 <= '1';
			out105 <= '1';
			out283 <= '1';
		end if;

		if state_cur(165) = '1' then
			-- Next state
			state_next(166) <= '1';
			-- Next values for buffered outputs
			out273_bufn <= '1';
			out343_bufn <= '1';
			out281_bufn <= '1';
			out181_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(166) = '1' then
			-- Next state
			state_next(215) <= '1';
			-- Next values for buffered outputs
			out562_bufn <= '1';
			out342_bufn <= '1';
			out284_bufn <= '1';
			out404_bufn <= '1';
			-- Assignment of non-buffered outputs
			out467 <= '1';
			out142 <= '1';
			out283 <= '1';
		end if;

		if state_cur(167) = '1' then
			if rtmcmp167 = '1' then
				-- Next state
				state_next(164) <= '1';
				-- Next values for buffered outputs
				out409_bufn <= '1';
				out351_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out130 <= '1';
				out101 <= '1';
				out112 <= '1';
				out142 <= '1';
				out99 <= '1';
				out54 <= '1';
				out135 <= '1';
				out123 <= '1';
				out114 <= '1';
				out286 <= '1';
			else  -- Stay in the current state
				state_next(167) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out475_bufn <= '1';
				out257_bufn <= '1';
				out472_bufn <= '1';
				out451_bufn <= '1';
				out468_bufn <= '1';
				out327_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out469 <= '1';
		end if;

		if state_cur(168) = '1' then
			-- Next state
			state_next(132) <= '1';
			-- Next values for buffered outputs
			out357_bufn <= '1';
			out428_bufn <= '1';
			out327_bufn <= '1';
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out283 <= '1';
		end if;

		if state_cur(169) = '1' then
			-- Next state
			state_next(225) <= '1';
			-- Next values for buffered outputs
			out554_bufn <= '1';
			out284_bufn <= '1';
			out333_bufn <= '1';
			-- Assignment of non-buffered outputs
			out137 <= '1';
			out135 <= '1';
			out484 <= '1';
			out283 <= '1';
		end if;

		if state_cur(170) = '1' then
			-- Next state
			state_next(152) <= '1';
			-- Next values for buffered outputs
			out353_bufn <= '1';
			out284_bufn <= '1';
			out138_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(171) = '1' then
			-- Next state
			state_next(167) <= '1';
			-- Next values for buffered outputs
			out475_bufn <= '1';
			out257_bufn <= '1';
			out472_bufn <= '1';
			out451_bufn <= '1';
			out468_bufn <= '1';
			out327_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(172) = '1' then
			-- Next state
			state_next(187) <= '1';
			-- Next values for buffered outputs
			out521_bufn <= '1';
			out284_bufn <= '1';
			out150_bufn <= '1';
			-- Assignment of non-buffered outputs
			out137 <= '1';
			out135 <= '1';
			out488 <= '1';
			out286 <= '1';
		end if;

		if state_cur(173) = '1' then
			-- Next state
			state_next(84) <= '1';
			-- Next values for buffered outputs
			out293_bufn <= '1';
			out281_bufn <= '1';
			out174_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(174) = '1' then
			if rtmcmp174 = '1' then
				-- Next state
				state_next(171) <= '1';
				-- Next values for buffered outputs
				out438_bufn <= '1';
				out324_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out125 <= '1';
				out137 <= '1';
				out116 <= '1';
				out56 <= '1';
				out283 <= '1';
			else  -- Stay in the current state
				state_next(174) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out229_bufn <= '1';
				out357_bufn <= '1';
				out407_bufn <= '1';
				out314_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out491 <= '1';
		end if;

		if state_cur(175) = '1' then
			-- Next state
			state_next(174) <= '1';
			-- Next values for buffered outputs
			out229_bufn <= '1';
			out357_bufn <= '1';
			out407_bufn <= '1';
			out314_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(176) = '1' then
			-- Next state
			state_next(175) <= '1';
			-- Next values for buffered outputs
			out495_bufn <= '1';
			out291_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(177) = '1' then
			-- Next state
			state_next(176) <= '1';
			-- Next values for buffered outputs
			out437_bufn <= '1';
			out289_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(178) = '1' then
			-- Next state
			state_next(145) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out103 <= '1';
			out105 <= '1';
			out99 <= '1';
			out101 <= '1';
		end if;

		if state_cur(179) = '1' then
			-- Next state
			state_next(177) <= '1';
			-- Next values for buffered outputs
			out496_bufn <= '1';
			out287_bufn <= '1';
			-- Assignment of non-buffered outputs
			out58 <= '1';
			out118 <= '1';
			out498 <= '1';
			out46 <= '1';
			out283 <= '1';
		end if;

		if state_cur(180) = '1' then
			-- Next state
			state_next(179) <= '1';
			-- Next values for buffered outputs
			out57_bufn <= '1';
			out497_bufn <= '1';
			out436_bufn <= '1';
			out294_bufn <= '1';
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out60 <= '1';
			out103 <= '1';
			out105 <= '1';
			out283 <= '1';
		end if;

		if state_cur(181) = '1' then
			if rtmcmp181 = '1' then
				-- Next state
				state_next(180) <= '1';
				-- Next values for buffered outputs
				out499_bufn <= '1';
				out351_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out130 <= '1';
				out101 <= '1';
				out112 <= '1';
				out142 <= '1';
				out99 <= '1';
				out54 <= '1';
				out135 <= '1';
				out123 <= '1';
				out114 <= '1';
				out286 <= '1';
			else  -- Stay in the current state
				state_next(181) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out260_bufn <= '1';
				out500_bufn <= '1';
				out435_bufn <= '1';
				out395_bufn <= '1';
				out327_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out501 <= '1';
		end if;

		if state_cur(182) = '1' then
			-- Next state
			state_next(181) <= '1';
			-- Next values for buffered outputs
			out260_bufn <= '1';
			out500_bufn <= '1';
			out435_bufn <= '1';
			out395_bufn <= '1';
			out327_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(183) = '1' then
			if rtmcmp183 = '1' then
				-- Next state
				state_next(182) <= '1';
				-- Next values for buffered outputs
				out457_bufn <= '1';
				out324_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out125 <= '1';
				out137 <= '1';
				out116 <= '1';
				out56 <= '1';
				out283 <= '1';
			else  -- Stay in the current state
				state_next(183) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out472_bufn <= '1';
				out401_bufn <= '1';
				out512_bufn <= '1';
				out314_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out513 <= '1';
		end if;

		if state_cur(184) = '1' then
			-- Next state
			state_next(183) <= '1';
			-- Next values for buffered outputs
			out472_bufn <= '1';
			out401_bufn <= '1';
			out512_bufn <= '1';
			out314_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(185) = '1' then
			-- Next state
			state_next(92) <= '1';
			-- Next values for buffered outputs
			out323_bufn <= '1';
			out284_bufn <= '1';
			out217_bufn <= '1';
			-- Assignment of non-buffered outputs
			out105 <= '1';
			out101 <= '1';
			out283 <= '1';
		end if;

		if state_cur(186) = '1' then
			-- Next state
			state_next(107) <= '1';
			-- Next values for buffered outputs
			out366_bufn <= '1';
			out315_bufn <= '1';
			out281_bufn <= '1';
			out183_bufn <= '1';
			-- Assignment of non-buffered outputs
			out142 <= '1';
			out519 <= '1';
			out286 <= '1';
		end if;

		if state_cur(187) = '1' then
			-- Next state
			state_next(185) <= '1';
			-- Next values for buffered outputs
			out290_bufn <= '1';
			out281_bufn <= '1';
			out248_bufn <= '1';
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out118 <= '1';
			out116 <= '1';
			out114 <= '1';
			out130 <= '1';
			out522 <= '1';
			out286 <= '1';
		end if;

		if state_cur(188) = '1' then
			-- Next state
			state_next(184) <= '1';
			-- Next values for buffered outputs
			out517_bufn <= '1';
			out291_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(189) = '1' then
			-- Next state
			state_next(190) <= '1';
			-- Next values for buffered outputs
			out526_bufn <= '1';
			out284_bufn <= '1';
			out213_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(190) = '1' then
			-- Next state
			state_next(173) <= '1';
			-- Next values for buffered outputs
			out468_bufn <= '1';
			out284_bufn <= '1';
			out143_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(191) = '1' then
			-- Next state
			state_next(188) <= '1';
			-- Next values for buffered outputs
			out524_bufn <= '1';
			out289_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(192) = '1' then
			-- Next state
			state_next(191) <= '1';
			-- Next values for buffered outputs
			out487_bufn <= '1';
			out287_bufn <= '1';
			-- Assignment of non-buffered outputs
			out58 <= '1';
			out118 <= '1';
			out527 <= '1';
			out44 <= '1';
			out283 <= '1';
		end if;

		if state_cur(193) = '1' then
			-- Next state
			state_next(192) <= '1';
			-- Next values for buffered outputs
			out57_bufn <= '1';
			out312_bufn <= '1';
			out433_bufn <= '1';
			out294_bufn <= '1';
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out60 <= '1';
			out103 <= '1';
			out105 <= '1';
			out283 <= '1';
		end if;

		if state_cur(194) = '1' then
			if rtmcmp194 = '1' then
				-- Next state
				state_next(193) <= '1';
				-- Next values for buffered outputs
				out351_bufn <= '1';
				out313_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out130 <= '1';
				out101 <= '1';
				out112 <= '1';
				out142 <= '1';
				out99 <= '1';
				out54 <= '1';
				out123 <= '1';
				out135 <= '1';
				out114 <= '1';
				out286 <= '1';
			else  -- Stay in the current state
				state_next(194) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out263_bufn <= '1';
				out531_bufn <= '1';
				out497_bufn <= '1';
				out521_bufn <= '1';
				out327_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out528 <= '1';
		end if;

		if state_cur(195) = '1' then
			-- Next state
			state_next(194) <= '1';
			-- Next values for buffered outputs
			out263_bufn <= '1';
			out531_bufn <= '1';
			out497_bufn <= '1';
			out521_bufn <= '1';
			out327_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(196) = '1' then
			-- Next state
			state_next(221) <= '1';
			-- Next values for buffered outputs
			out281_bufn <= '1';
			-- Assignment of non-buffered outputs
			out130 <= '1';
			out540 <= '1';
			out286 <= '1';
		end if;

		if state_cur(197) = '1' then
			if rtmcmp197 = '1' then
				-- Next state
				state_next(195) <= '1';
				-- Next values for buffered outputs
				out394_bufn <= '1';
				out324_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out137 <= '1';
				out125 <= '1';
				out116 <= '1';
				out56 <= '1';
				out283 <= '1';
			else  -- Stay in the current state
				state_next(197) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out500_bufn <= '1';
				out435_bufn <= '1';
				out314_bufn <= '1';
				out293_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out542 <= '1';
		end if;

		if state_cur(198) = '1' then
			-- Next state
			state_next(197) <= '1';
			-- Next values for buffered outputs
			out500_bufn <= '1';
			out435_bufn <= '1';
			out314_bufn <= '1';
			out293_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(199) = '1' then
			-- Next state
			state_next(198) <= '1';
			-- Next values for buffered outputs
			out326_bufn <= '1';
			out291_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(200) = '1' then
			-- Next state
			state_next(199) <= '1';
			-- Next values for buffered outputs
			out341_bufn <= '1';
			out289_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(201) = '1' then
			-- Next state
			state_next(200) <= '1';
			-- Next values for buffered outputs
			out287_bufn <= '1';
			out285_bufn <= '1';
			-- Assignment of non-buffered outputs
			out58 <= '1';
			out118 <= '1';
			out544 <= '1';
			out42 <= '1';
			out283 <= '1';
		end if;

		if state_cur(202) = '1' then
			-- Next state
			state_next(201) <= '1';
			-- Next values for buffered outputs
			out57_bufn <= '1';
			out318_bufn <= '1';
			out322_bufn <= '1';
			out294_bufn <= '1';
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out60 <= '1';
			out103 <= '1';
			out105 <= '1';
			out283 <= '1';
		end if;

		if state_cur(203) = '1' then
			if rtmcmp203 = '1' then
				-- Next state
				state_next(202) <= '1';
				-- Next values for buffered outputs
				out483_bufn <= '1';
				out351_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out130 <= '1';
				out101 <= '1';
				out142 <= '1';
				out112 <= '1';
				out99 <= '1';
				out54 <= '1';
				out123 <= '1';
				out135 <= '1';
				out114 <= '1';
				out286 <= '1';
			else  -- Stay in the current state
				state_next(203) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out393_bufn <= '1';
				out346_bufn <= '1';
				out344_bufn <= '1';
				out312_bufn <= '1';
				out518_bufn <= '1';
				out327_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out545 <= '1';
		end if;

		if state_cur(204) = '1' then
			-- Next state
			state_next(203) <= '1';
			-- Next values for buffered outputs
			out393_bufn <= '1';
			out346_bufn <= '1';
			out344_bufn <= '1';
			out312_bufn <= '1';
			out518_bufn <= '1';
			out327_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(205) = '1' then
			if rtmcmp205 = '1' then
				-- Next state
				state_next(204) <= '1';
				-- Next values for buffered outputs
				out554_bufn <= '1';
				out324_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out137 <= '1';
				out125 <= '1';
				out116 <= '1';
				out56 <= '1';
				out283 <= '1';
			else  -- Stay in the current state
				state_next(205) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out531_bufn <= '1';
				out426_bufn <= '1';
				out461_bufn <= '1';
				out314_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out555 <= '1';
		end if;

		if state_cur(206) = '1' then
			-- Next state
			state_next(205) <= '1';
			-- Next values for buffered outputs
			out531_bufn <= '1';
			out426_bufn <= '1';
			out461_bufn <= '1';
			out314_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(207) = '1' then
			-- Next state
			state_next(206) <= '1';
			-- Next values for buffered outputs
			out526_bufn <= '1';
			out291_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(208) = '1' then
			-- Next state
			state_next(207) <= '1';
			-- Next values for buffered outputs
			out525_bufn <= '1';
			out289_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(209) = '1' then
			-- Next state
			state_next(208) <= '1';
			-- Next values for buffered outputs
			out466_bufn <= '1';
			out287_bufn <= '1';
			-- Assignment of non-buffered outputs
			out58 <= '1';
			out118 <= '1';
			out559 <= '1';
			out40 <= '1';
			out283 <= '1';
		end if;

		if state_cur(210) = '1' then
			-- Next state
			state_next(209) <= '1';
			-- Next values for buffered outputs
			out57_bufn <= '1';
			out417_bufn <= '1';
			out294_bufn <= '1';
			out282_bufn <= '1';
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out60 <= '1';
			out103 <= '1';
			out105 <= '1';
			out283 <= '1';
		end if;

		if state_cur(211) = '1' then
			-- Next state
			state_next(224) <= '1';
			-- Next values for buffered outputs
			out459_bufn <= '1';
			out284_bufn <= '1';
			out201_bufn <= '1';
			-- Assignment of non-buffered outputs
			out560 <= '1';
			out286 <= '1';
		end if;

		if state_cur(212) = '1' then
			-- Next state
			state_next(147) <= '1';
			-- Next values for buffered outputs
			out49_bufn <= '1';
			-- Assignment of non-buffered outputs
			out60 <= '1';
			out561 <= '1';
			out58 <= '1';
			out56 <= '1';
			out54 <= '1';
		end if;

		if state_cur(213) = '1' then
			-- Next state
			state_next(134) <= '1';
			-- Next values for buffered outputs
			out433_bufn <= '1';
			out281_bufn <= '1';
			out426_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(214) = '1' then
			-- Next state
			state_next(140) <= '1';
			-- Next values for buffered outputs
			out351_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(215) = '1' then
			if rtmcmp215 = '1' then
				-- Next state
				state_next(127) <= '1';
				-- Next values for buffered outputs
				out404_bufn <= '1';
				out418_bufn <= '1';
				out281_bufn <= '1';
				out417_bufn <= '1';
				-- Last cycle of current state: assignment of non-buffered outputs
				out125 <= '1';
				out123 <= '1';
				out286 <= '1';
			else  -- Stay in the current state
				state_next(215) <= '1';
				rtmcounter0_next <= rtmcounter0 + 1;
				-- Maintain buffered outputs
				out562_bufn <= '1';
				out342_bufn <= '1';
				out284_bufn <= '1';
				out404_bufn <= '1';
			end if;
			-- Assignment of non-buffered outputs;
				out563 <= '1';
		end if;

		if state_cur(216) = '1' then
			-- Next state
			state_next(214) <= '1';
			-- Next values for buffered outputs
			out482_bufn <= '1';
			out481_bufn <= '1';
			out357_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(217) = '1' then
			-- Next state
			state_next(216) <= '1';
			-- Next values for buffered outputs
			out444_bufn <= '1';
			out281_bufn <= '1';
			out354_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(218) = '1' then
			-- Next state
			state_next(217) <= '1';
			-- Next values for buffered outputs
			out566_bufn <= '1';
			out281_bufn <= '1';
			out229_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(219) = '1' then
			-- Next state
			state_next(218) <= '1';
			-- Next values for buffered outputs
			out440_bufn <= '1';
			out281_bufn <= '1';
			out162_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(220) = '1' then
			-- Next state
			state_next(219) <= '1';
			-- Next values for buffered outputs
			out349_bufn <= '1';
			out284_bufn <= '1';
			out257_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(221) = '1' then
			-- Next state
			state_next(223) <= '1';
			-- Next values for buffered outputs
			out325_bufn <= '1';
			out284_bufn <= '1';
			out366_bufn <= '1';
			-- Assignment of non-buffered outputs
			out112 <= '1';
			out567 <= '1';
			out283 <= '1';
		end if;

		if state_cur(222) = '1' then
			-- Next state
			state_next(220) <= '1';
			-- Next values for buffered outputs
			out464_bufn <= '1';
			out281_bufn <= '1';
			out451_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(223) = '1' then
			-- Next state
			state_next(161) <= '1';
			-- Next values for buffered outputs
			out57_bufn <= '1';
			out414_bufn <= '1';
			out446_bufn <= '1';
			-- Assignment of non-buffered outputs
			out105 <= '1';
			out103 <= '1';
			out101 <= '1';
			out99 <= '1';
			out286 <= '1';
		end if;

		if state_cur(224) = '1' then
			-- Next state
			state_next(222) <= '1';
			-- Next values for buffered outputs
			out460_bufn <= '1';
			out281_bufn <= '1';
			out232_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(225) = '1' then
			-- Next state
			state_next(79) <= '1';
			-- Next values for buffered outputs
			out282_bufn <= '1';
			out281_bufn <= '1';
			out280_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(226) = '1' then
			-- Next state
			state_next(122) <= '1';
			-- Next values for buffered outputs
			out111_bufn <= '1';
			out410_bufn <= '1';
			-- Assignment of non-buffered outputs
			out52 <= '1';
			out21 <= '1';
			out125 <= '1';
			out123 <= '1';
			out570 <= '1';
			out412 <= '1';
		end if;

		if state_cur(227) = '1' then
			-- Next state
			state_next(116) <= '1';
			-- Next values for buffered outputs
			out400_bufn <= '1';
			out284_bufn <= '1';
			out131_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(228) = '1' then
			-- Next state
			state_next(136) <= '1';
			-- Next values for buffered outputs
			out428_bufn <= '1';
			out284_bufn <= '1';
			out126_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(229) = '1' then
			-- Next state
			state_next(138) <= '1';
			-- Next values for buffered outputs
			out437_bufn <= '1';
			out281_bufn <= '1';
			out235_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(230) = '1' then
			-- Next state
			state_next(231) <= '1';
			-- Next values for buffered outputs
			out499_bufn <= '1';
			out281_bufn <= '1';
			out497_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(231) = '1' then
			-- Next state
			state_next(155) <= '1';
			-- Next values for buffered outputs
			out457_bufn <= '1';
			out284_bufn <= '1';
			out364_bufn <= '1';
			-- Assignment of non-buffered outputs
			out283 <= '1';
		end if;

		if state_cur(232) = '1' then
			-- Next state
			state_next(213) <= '1';
			-- Next values for buffered outputs
			out524_bufn <= '1';
			out281_bufn <= '1';
			out238_bufn <= '1';
			-- Assignment of non-buffered outputs
			out286 <= '1';
		end if;

		if state_cur(233) = '1' then
			-- Next state
			state_next(141) <= '1';
			-- Next values for buffered outputs
			out440_bufn <= '1';
			out314_bufn <= '1';
			-- Assignment of non-buffered outputs
			out118 <= '1';
			out283 <= '1';
		end if;

		if state_cur(234) = '1' then
			-- Next state
			state_next(129) <= '1';
			-- Next values for buffered outputs
			out346_bufn <= '1';
			out31_bufn <= '1';
			out410_bufn <= '1';
			-- Assignment of non-buffered outputs
			out42 <= '1';
			out21 <= '1';
			out572 <= '1';
			out412 <= '1';
		end if;

		if state_cur(235) = '1' then
			-- Next state
			state_next(131) <= '1';
			-- Next values for buffered outputs
			-- Assignment of non-buffered outputs
			out120 <= '1';
			out118 <= '1';
			out116 <= '1';
			out114 <= '1';
			out112 <= '1';
			out575 <= '1';
			out363 <= '1';
		end if;

		if state_cur(236) = '1' then
			-- Next state
			state_next(234) <= '1';
			-- Next values for buffered outputs
			out280_bufn <= '1';
			out410_bufn <= '1';
			-- Assignment of non-buffered outputs
			out577 <= '1';
			out40 <= '1';
			out21 <= '1';
			out412 <= '1';
		end if;

		if state_cur(237) = '1' then
			-- Next state
			state_next(235) <= '1';
			-- Next values for buffered outputs
			out111_bufn <= '1';
			out361_bufn <= '1';
			-- Assignment of non-buffered outputs
			out52 <= '1';
			out21 <= '1';
			out125 <= '1';
			out123 <= '1';
			out578 <= '1';
			out363 <= '1';
		end if;

		if state_cur(238) = '1' then
			-- Next state
			state_next(236) <= '1';
			-- Next values for buffered outputs
			out562_bufn <= '1';
			out35_bufn <= '1';
			out410_bufn <= '1';
			-- Assignment of non-buffered outputs
			out580 <= '1';
			out38 <= '1';
			out21 <= '1';
		end if;

		if state_cur(239) = '1' then
			-- Next state
			state_next(238) <= '1';
			-- Next values for buffered outputs
			out446_bufn <= '1';
			out36_bufn <= '1';
			-- Assignment of non-buffered outputs
			out50 <= '1';
			out46 <= '1';
			out52 <= '1';
			out48 <= '1';
			out44 <= '1';
			out42 <= '1';
			out40 <= '1';
			out38 <= '1';
		end if;

		if state_cur(240) = '1' then
			-- Next state
			state_next(165) <= '1';
			-- Next values for buffered outputs
			out466_bufn <= '1';
			out284_bufn <= '1';
			out273_bufn <= '1';
			-- Assignment of non-buffered outputs
			out581 <= '1';
			out130 <= '1';
			out283 <= '1';
		end if;

		-- Reset input
		if reset = '1' then
			-- Set the reset state
			state_next <= (7 => '1', others => '0');
			-- Note: Resetting all buffers for outputs here is not necessary.
			-- It would cost hardware. They will be reset at the next clock front.
			-- Retiming: counters
			rtmcounter0_next <= (others => '0');
			-- Reset state: set the buffered outputs
		end if;

	end process;

	-- Assignment of buffered outputs

	out122 <= out122_buf;
	out36 <= out36_buf;
	out49 <= out49_buf;
	out35 <= out35_buf;
	out27 <= out27_buf;
	out16 <= out16_buf;
	out25 <= out25_buf;
	out20 <= out20_buf;
	out57 <= out57_buf;
	out23 <= out23_buf;
	out136 <= out136_buf;
	out0 <= out0_buf;
	out134 <= out134_buf;
	out13 <= out13_buf;
	out131 <= out131_buf;
	out129 <= out129_buf;
	out111 <= out111_buf;
	out31 <= out31_buf;
	out126 <= out126_buf;
	out106 <= out106_buf;
	out124 <= out124_buf;
	out138 <= out138_buf;
	out141 <= out141_buf;
	out143 <= out143_buf;
	out146 <= out146_buf;
	out150 <= out150_buf;
	out153 <= out153_buf;
	out155 <= out155_buf;
	out158 <= out158_buf;
	out162 <= out162_buf;
	out165 <= out165_buf;
	out168 <= out168_buf;
	out171 <= out171_buf;
	out174 <= out174_buf;
	out178 <= out178_buf;
	out181 <= out181_buf;
	out183 <= out183_buf;
	out197 <= out197_buf;
	out201 <= out201_buf;
	out204 <= out204_buf;
	out207 <= out207_buf;
	out210 <= out210_buf;
	out213 <= out213_buf;
	out217 <= out217_buf;
	out220 <= out220_buf;
	out222 <= out222_buf;
	out225 <= out225_buf;
	out229 <= out229_buf;
	out232 <= out232_buf;
	out235 <= out235_buf;
	out238 <= out238_buf;
	out241 <= out241_buf;
	out245 <= out245_buf;
	out248 <= out248_buf;
	out250 <= out250_buf;
	out253 <= out253_buf;
	out257 <= out257_buf;
	out260 <= out260_buf;
	out263 <= out263_buf;
	out266 <= out266_buf;
	out269 <= out269_buf;
	out273 <= out273_buf;
	out276 <= out276_buf;
	out278 <= out278_buf;
	out280 <= out280_buf;
	out281 <= out281_buf;
	out282 <= out282_buf;
	out284 <= out284_buf;
	out285 <= out285_buf;
	out287 <= out287_buf;
	out288 <= out288_buf;
	out289 <= out289_buf;
	out290 <= out290_buf;
	out291 <= out291_buf;
	out292 <= out292_buf;
	out293 <= out293_buf;
	out294 <= out294_buf;
	out295 <= out295_buf;
	out296 <= out296_buf;
	out312 <= out312_buf;
	out313 <= out313_buf;
	out314 <= out314_buf;
	out315 <= out315_buf;
	out318 <= out318_buf;
	out322 <= out322_buf;
	out323 <= out323_buf;
	out324 <= out324_buf;
	out325 <= out325_buf;
	out326 <= out326_buf;
	out327 <= out327_buf;
	out328 <= out328_buf;
	out333 <= out333_buf;
	out341 <= out341_buf;
	out342 <= out342_buf;
	out343 <= out343_buf;
	out344 <= out344_buf;
	out346 <= out346_buf;
	out349 <= out349_buf;
	out351 <= out351_buf;
	out352 <= out352_buf;
	out353 <= out353_buf;
	out354 <= out354_buf;
	out357 <= out357_buf;
	out361 <= out361_buf;
	out364 <= out364_buf;
	out366 <= out366_buf;
	out371 <= out371_buf;
	out393 <= out393_buf;
	out394 <= out394_buf;
	out395 <= out395_buf;
	out400 <= out400_buf;
	out401 <= out401_buf;
	out404 <= out404_buf;
	out407 <= out407_buf;
	out408 <= out408_buf;
	out409 <= out409_buf;
	out410 <= out410_buf;
	out413 <= out413_buf;
	out414 <= out414_buf;
	out417 <= out417_buf;
	out418 <= out418_buf;
	out422 <= out422_buf;
	out426 <= out426_buf;
	out428 <= out428_buf;
	out431 <= out431_buf;
	out433 <= out433_buf;
	out434 <= out434_buf;
	out435 <= out435_buf;
	out436 <= out436_buf;
	out437 <= out437_buf;
	out438 <= out438_buf;
	out440 <= out440_buf;
	out444 <= out444_buf;
	out446 <= out446_buf;
	out451 <= out451_buf;
	out457 <= out457_buf;
	out458 <= out458_buf;
	out459 <= out459_buf;
	out460 <= out460_buf;
	out461 <= out461_buf;
	out463 <= out463_buf;
	out464 <= out464_buf;
	out466 <= out466_buf;
	out468 <= out468_buf;
	out472 <= out472_buf;
	out475 <= out475_buf;
	out481 <= out481_buf;
	out482 <= out482_buf;
	out483 <= out483_buf;
	out487 <= out487_buf;
	out495 <= out495_buf;
	out496 <= out496_buf;
	out497 <= out497_buf;
	out499 <= out499_buf;
	out500 <= out500_buf;
	out512 <= out512_buf;
	out517 <= out517_buf;
	out518 <= out518_buf;
	out521 <= out521_buf;
	out524 <= out524_buf;
	out525 <= out525_buf;
	out526 <= out526_buf;
	out531 <= out531_buf;
	out554 <= out554_buf;
	out562 <= out562_buf;
	out566 <= out566_buf;

	-- Retiming: the comparators

	rtmcmp90 <= '1' when state_cur(90) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp95 <= '1' when state_cur(95) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp98 <= '1' when state_cur(98) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp104 <= '1' when state_cur(104) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp148 <= '1' when state_cur(148) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp167 <= '1' when state_cur(167) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp174 <= '1' when state_cur(174) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp181 <= '1' when state_cur(181) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp183 <= '1' when state_cur(183) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp194 <= '1' when state_cur(194) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp197 <= '1' when state_cur(197) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp203 <= '1' when state_cur(203) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp205 <= '1' when state_cur(205) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp215 <= '1' when state_cur(215) = '1' and rtmcounter0 = 1 else '0';

end architecture;

