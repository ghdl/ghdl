
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2853.vhd,v 1.2 2001-10-26 16:29:49 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c13s10b00x00p02n01i02853ent IS
END c13s10b00x00p02n01i02853ent;

ARCHITECTURE c13s10b00x00p02n01i02853arch OF c13s10b00x00p02n01i02853ent IS

BEGIN
  TESTING: PROCESS
    subtype   BYTE is BIT_VECTOR (0 to 7);
    variable   b1 : BYTE;
    variable    b2 : BYTE;
  BEGIN
    b1 := BYTE'(0 | 1 | 2 | 3 | 4 | 5 | 6 | 7 => '1');
    b2 := BYTE'(0 ! 1 ! 2 ! 3 ! 4 ! 5 ! 6 ! 7 => '1');
    assert NOT( b1=b2 )
      report "***PASSED TEST: c13s10b00x00p02n01i02853"
      severity NOTE;
    assert ( b1=b2 )
      report "***FAILED TEST: c13s10b00x00p02n01i02853 - "
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c13s10b00x00p02n01i02853arch;
