entity mwe is
end entity;

architecture test of mwe is
    signal b : bit;
begin
end architecture;
