entity tb is
end tb;

architecture behavioral of tb is
  function A(v : integer) return i000'er is
  begin
  end;
begin
end behavioral;

