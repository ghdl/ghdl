
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc179.vhd,v 1.2 2001-10-26 16:29:43 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c04s04b00x00p02n01i00179ent IS
  attribute attr : INTEGER;
END c04s04b00x00p02n01i00179ent;

ARCHITECTURE c04s04b00x00p02n01i00179arch OF c04s04b00x00p02n01i00179ent IS
  constant    C : INTEGER    := 1;
  attribute    attr of C : CONSTANT       is 40;
  constant    D : INTEGER    := C'attr;
BEGIN
  TESTING: PROCESS
  BEGIN
    wait for 5 ns;
    assert NOT( C = 1 and D = 40 )
      report "***PASSED TEST: c04s04b00x00p02n01i00179"
      severity NOTE;
    assert ( C = 1 and D = 40 )
      report "***FAILED TEST: c04s04b00x00p02n01i00179 - User-defined attribute test failed."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c04s04b00x00p02n01i00179arch;
