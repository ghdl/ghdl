
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc318.vhd,v 1.2 2001-10-26 16:29:52 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s02b01x00p03n01i00318ent IS
END c03s02b01x00p03n01i00318ent;

ARCHITECTURE c03s02b01x00p03n01i00318arch OF c03s02b01x00p03n01i00318ent IS
  type MVL is ('0', '1', 'Z') ;
  type MVL_vector is array (0 to 63)of MVL;
BEGIN
  TESTING: PROCESS
    variable k : MVL_vector;
  BEGIN
    k(5) := 'Z';
    assert NOT(k(5)='Z')
      report "***PASSED TEST: c03s02b01x00p03n01i00318"
      severity NOTE;
    assert (k(5)='Z')
      report "***FAILED TEST: c03s02b01x00p03n01i00318 - In the unconstrained array definition, the reserved word array has been followed by a list of index subtype definitions enclosed with parentheses and the reserved word of."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s02b01x00p03n01i00318arch;
