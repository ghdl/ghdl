library ieee;
use ieee.std_logic_arith.all;

entity tb is
end tb;
