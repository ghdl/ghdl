entity ent is
end entity;

architecture a of ent is
begin
 -- Comment added.
end architecture;
