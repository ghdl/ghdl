
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc3014.vhd,v 1.2 2001-10-26 16:30:24 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

package c11s01b00x00p08n03i03014ent is
  procedure test;
end c11s01b00x00p08n03i03014ent;

package body c11s01b00x00p08n03i03014ent is
  procedure test  is
  begin
    assert false
      report "Duplicate primary unit name allowed in same library -- test fails."
      severity note ;
  end test;
end c11s01b00x00p08n03i03014ent;

use work.c11s01b00x00p08n03i03014ent.all;
ENTITY c11s01b00x00p08n03i03014ent IS
END c11s01b00x00p08n03i03014ent;

ARCHITECTURE c11s01b00x00p08n03i03014arch OF c11s01b00x00p08n03i03014ent IS

BEGIN
  c11s01b00x00p08n03i03014ent.test;

  TESTING: PROCESS
  BEGIN
    assert FALSE
      report "***FAILED TEST: c11s01b00x00p08n03i03014d - Duplicate primary unit name is not allowed in same library."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c11s01b00x00p08n03i03014arch;
