
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1322.vhd,v 1.2 2001-10-26 16:29:40 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c08s04b00x00p09n04i01322ent IS
END c08s04b00x00p09n04i01322ent;

ARCHITECTURE c08s04b00x00p09n04i01322arch OF c08s04b00x00p09n04i01322ent IS
  signal S1 : BIT := '1';
  signal S2 : BIT := '1';
BEGIN
  S1 <= transport '0' after 5 ns,
        '1' after 10 ns;
  S2 <= S1 after 15 ns;
  TESTING: PROCESS(S2)
  BEGIN
    assert NOT( S2 = '1' )
      report "***PASSED TEST: c08s04b00x00p09n04i01322"
      severity NOTE;
    assert ( S2 = '1' )
      report "***FAILED TEST: c08s04b00x00p09n04i01322 - A pulse whose duration is shorter than the switching time of the circuit is not transmitted."
      severity ERROR;
  END PROCESS TESTING;

END c08s04b00x00p09n04i01322arch;
