
-- Copyright (C) 2002 Morgan Kaufmann Publishers, Inc

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

library ieee_proposed;  use ieee_proposed.electrical_systems.all;
                        
entity mixer is
  port ( terminal inputs : electrical_vector(1 to 8);
         terminal output : electrical );
end entity mixer;

----------------------------------------------------------------

architecture weighted of mixer is
  
  quantity v_in across inputs;
  quantity v_out across i_out through output;
  constant gains : real_vector(1 to 8)
    := ( 0.01, 0.04, 0.15, 0.30, 0.03, 0.15, 0.04, 0.01 );
  
begin
  
  apply_weights : procedural is
    variable sum : real := 0.0;
  begin
    for index in v_in'range loop
      sum := sum + v_in(index) * gains(index);
    end loop;
    v_out := sum;
  end procedural apply_weights;
        
end architecture weighted;
