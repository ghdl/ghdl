
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc927.vhd,v 1.2 2001-10-26 16:30:02 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

package c10s04b00x00p01n01i00927pkg is
  type work is array(0 to 7) of BIT;
end c10s04b00x00p01n01i00927pkg;

use  work.c10s04b00x00p01n01i00927pkg.all;
ENTITY c10s04b00x00p01n01i00927ent IS
  port (P : in  bit);
END c10s04b00x00p01n01i00927ent;

ARCHITECTURE c10s04b00x00p01n01i00927arch OF c10s04b00x00p01n01i00927ent IS
  use  work.c10s04b00x00p01n01i00927pkg;
BEGIN
  TESTING: PROCESS(P)
    -- This succeeds because type work is defined in package c10s04b00x00p01n01i00927pkg,
    -- there is no conflict with library "work"
    variable doit : c10s04b00x00p01n01i00927pkg.work ;  -- No_failure_here
  BEGIN
    assert NOT(doit="00000000") 
      report "***PASSED TEST: c10s04b00x00p01n01i00927"
      severity NOTE;
    assert (doit="00000000") 
      report "***FAILED TEST: c10s04b00x00p01n01i00927 - Use clause do not make that declaration visible." 
      severity ERROR;
  END PROCESS TESTING;

END c10s04b00x00p01n01i00927arch;
