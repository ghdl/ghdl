entity function()return n(of