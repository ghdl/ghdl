
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc265.vhd,v 1.2 2001-10-26 16:29:49 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s01b03x00p02n01i00265ent IS
END c03s01b03x00p02n01i00265ent;

ARCHITECTURE c03s01b03x00p02n01i00265arch OF c03s01b03x00p02n01i00265ent IS
  type J is           -- physical type decl
    range 0 to 1000
    units
      A;
      B = 10 A;
      C = 10 B;
      D = 10 C;
    end units;
  type J1 is access J;   -- Success_here
BEGIN
  TESTING: PROCESS
    variable k : J; 
  BEGIN
    k := 10 C;
    assert NOT( k=100 B )
      report "***PASSED TEST: c03s01b03x00p02n01i00265"
      severity NOTE;
    assert ( k=100 B)
      report "***FAILED TEST: c03s01b03x00p02n01i00265 - In the physical type definition, the range constraint is immediately followed by reserved word units."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s01b03x00p02n01i00265arch;
