package pkga is
  subtype word is bit_vector (31 downto 0);
end pkga;

