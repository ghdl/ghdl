entity tb is
end tb;

use work.pkg0.all;
use work.pkg1.all;
use work.pkg2.all;
use work.pkg3.all;
use work.pkg5.all;

architecture behav of tb is
begin
end behav;
