entity tb is
end;

architecture behav of tb is
begin
  assert 0!;
end behav;
