
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1127.vhd,v 1.2 2001-10-26 16:30:06 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c06s05b00x00p04n01i01127ent IS
END c06s05b00x00p04n01i01127ent;

ARCHITECTURE c06s05b00x00p04n01i01127arch OF c06s05b00x00p04n01i01127ent IS

  type idx is range 1 to 10;
  type aray1 is array (idx) of bit;
  type aray2 is array (idx range <>) of aray1;
BEGIN
  TESTING: PROCESS
    variable v2 : aray1;
    variable v3 : aray2(1 to 2);
  BEGIN
    v2 := v3(2 to 2)(1);             -- wrong index
    assert FALSE 
      report "***FAILED TEST: c06s05b00x00p04n01i01127 - Invalid index for slice." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c06s05b00x00p04n01i01127arch;
