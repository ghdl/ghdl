
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1149.vhd,v 1.2 2001-10-26 16:29:39 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c06s05b00x00p07n02i01149ent IS
END c06s05b00x00p07n02i01149ent;

ARCHITECTURE c06s05b00x00p07n02i01149arch OF c06s05b00x00p07n02i01149ent IS
  type    A is array (10 downto 1) of integer;
BEGIN
  TESTING: PROCESS
    variable var : A := (66,66,others=>6);
  BEGIN
    wait for 5 ns;
    assert NOT( var(1) = 6 )
      report "***PASSED TEST: c06s05b00x00p07n02i01149"
      severity NOTE;
    assert ( var(1) = 6 )
      report "***FAILED TEST: c06s05b00x00p07n02i01149 - A(N) is an element of the array A(decline) and has the corresponding element type."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c06s05b00x00p07n02i01149arch;
