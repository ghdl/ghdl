entity inter1 is
  port (variable a : boolean);
end inter1;
