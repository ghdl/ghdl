entity reserved2 is
end;

architecture behav of reserved2 is
  signal context : bit;
begin
  process
  begin
    wait;
  end process;
end behav;
