
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc30.vhd,v 1.2 2001-10-26 16:29:50 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c04s03b00x00p14n04i00030ent IS
END c04s03b00x00p14n04i00030ent;

ARCHITECTURE c04s03b00x00p14n04i00030arch OF c04s03b00x00p14n04i00030ent IS
  signal       M1 : BIT_VECTOR(0 to 7) ;
  constant    M2 : BIT := '1' ;
BEGIN
  TESTING: PROCESS
    variable   V1 : BIT; 
  BEGIN
    M1(3) <=    '1' after 10 ns;
    --- No_failure_here
    --- M1(3) is also a signal; so this signal
    --- assignment is possible.
    V1    :=    M2;   
    wait for 10 ns;
    assert NOT( M1(3)='1' and V1='1' )
      report "***PASSED TEST: c04s03b00x00p14n04i00030"
      severity NOTE;
    assert ( M1(3)='1' and V1='1' )
      report "***FAILED TEST:c04s03b00x00p14n04i00030 - Each subelement of that object is itself an object of the same class as the given object."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c04s03b00x00p14n04i00030arch;
