entity crash1 is
end crash1;

architecture behav of crash1 is
  signal samples: bit;
begin
  process
  begin
    bit'(samples));
  end process;
end behav;
