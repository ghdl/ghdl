package function is
if)n';