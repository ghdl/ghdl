
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2736.vhd,v 1.2 2001-10-26 16:29:49 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c13s06b00x00p01n01i02736ent IS
END c13s06b00x00p01n01i02736ent;

ARCHITECTURE c13s06b00x00p01n01i02736arch OF c13s06b00x00p01n01i02736ent IS

BEGIN
  TESTING: PROCESS
    variable S45 : STRING (1 to 44);
    variable S50 : STRING (1 to 50);
  BEGIN
    S45 := "ABCDEFGHIJKLMNOPQRSTUVWXYZ0123456789#&'()*+,";
    S50 := "-./:;<=>_| abcdefghijklmnopqrstuvwxyz!$%@?[\]^`{}~";
    wait for 5 ns;
    assert NOT(       S45 = "ABCDEFGHIJKLMNOPQRSTUVWXYZ0123456789#&'()*+,"
                      and S50 = "-./:;<=>_| abcdefghijklmnopqrstuvwxyz!$%@?[\]^`{}~")
      report "***PASSED TEST: c13s06b00x00p01n01i02736"
      severity NOTE;
    assert (       S45 = "ABCDEFGHIJKLMNOPQRSTUVWXYZ0123456789#&'()*+,"
                   and S50 = "-./:;<=>_| abcdefghijklmnopqrstuvwxyz!$%@?[\]^`{}~")
      report "***FAILED TEST: c13s06b00x00p01n01i02736 - String literal lexical test failed."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c13s06b00x00p01n01i02736arch;
