package p is
  type state_t is
    (
      s1,  --  For :s1:
      s2,
      s3  --  For :s3:
      );
end p;
