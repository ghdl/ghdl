entity libparen is
end libparen;

architecture behav of libparen is
  constant c : boolean := work(5);
begin
end behav;
