
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc162.vhd,v 1.2 2001-10-26 16:29:42 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

package c04s03b02x02p20n02i00162pkg is
  subtype string_v is string(1 to 32);
  CONSTANT null_string_v : string_v := (
    'A', 'B', 'C', 'D', 'E', 'F', 'G', 'H', 'I', 'J', 'K', 'L', 'M', 'N', 'O', 'P',
    'Q', 'R', 'S', 'T', 'U', 'V', 'W', 'X', 'Y', 'Z', 'a', 'b', 'c', 'd', 'e', 'f');
end c04s03b02x02p20n02i00162pkg;

ENTITY c04s03b02x02p20n02i00162ent IS
END c04s03b02x02p20n02i00162ent;

use work.c04s03b02x02p20n02i00162pkg.all;
ARCHITECTURE c04s03b02x02p20n02i00162arch OF c04s03b02x02p20n02i00162ent IS

BEGIN
  TESTING: PROCESS
    variable buf : string_v := null_string_v; 

    PROCEDURE sprintf
      (
        buff   : out string_v;
        str1   : in  string := null_string_v;
        str2   : in  string := null_string_v;
        str3   : in  string := null_string_v
        )
    is
      VARIABLE index : integer := 1;
    begin

      buff := null_string_v;

      for i in str1'range LOOP
        exit when str1(i) = ' ';
        buff (index) := str1 (i);
        index := index + 1;
      end LOOP;
      for i in str2'range LOOP
        exit when str2(i) = ' ';
        buff (index) := str2 (i);
        index := index + 1;
      end LOOP;
      for i in str3'range LOOP
        exit when str3(i) = ' ';
        buff (index) := str3 (i);
        index := index + 1;
      end LOOP;
    end sprintf;

  BEGIN
    sprintf ( buf,
              "VHDL ",
              "TECHNOLOGY ",
              "GROUP " );
    wait for 10 ns;

    assert NOT( buf(1  to 19) = "VHDLTECHNOLOGYGROUP"   and
                buf(20 to 32) = "TUVWXYZabcdef")
      report "***PASSED TEST: c04s03b02x02p20n02i00162"
      severity NOTE;
    assert ( buf(1  to 19) = "VHDLTECHNOLOGYGROUP"   and
             buf(20 to 32) = "TUVWXYZabcdef")
      report "***FAILED TEST: c04s03b02x02p20n02i00162- The value of the default expression is used as the actual expression in an implicit association element fot that interface element."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c04s03b02x02p20n02i00162arch;
