entity ent is
end entity;

architecture a of ent is
begin
  main : process
  begin
    report "Hello World";
    wait;
  end process;
end architecture;
