
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1975.vhd,v 1.2 2001-10-26 16:29:44 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c07s02b01x00p02n02i01975ent IS
  constant T:bit := '1';
  constant F:bit := '0';
END c07s02b01x00p02n02i01975ent;

ARCHITECTURE c07s02b01x00p02n02i01975arch OF c07s02b01x00p02n02i01975ent IS

BEGIN
  TESTING: PROCESS
    variable A1 : bit := T;
    variable A2 : bit := F;
  BEGIN
    assert NOT(    (A1 and A1) = '1'   and
                   (A1 and A2) = '0'   and
                   (A2 and A1) = '0'   and
                   (A2 and A2) = '0'   and
                   (A1 or A1) = '1'   and
                   (A1 or A2) = '1'   and
                   (A2 or A1) = '1'   and
                   (A2 or A2) = '0'   and
                   (A1 xor A1) = '0'   and
                   (A1 xor A2) = '1'   and
                   (A2 xor A1) = '1'   and
                   (A2 xor A2) = '0'   and
                   (A1 nand A1) = '0'   and
                   (A1 nand A2) = '1'   and
                   (A2 nand A1) = '1'   and
                   (A2 nand A2) = '1'   and
                   (A1 nor A1) = '0'   and
                   (A1 nor A2) = '0'   and
                   (A2 nor A1) = '0'   and
                   (A2 nor A2) = '1'   and
                   (not A1) = '0'      and
                   (not A2) = '1')
      report "***PASSED TEST: c07s02b01x00p02n02i01975"
      severity NOTE;
    assert (    (A1 and A1) = '1'   and
                (A1 and A2) = '0'   and
                (A2 and A1) = '0'   and
                (A2 and A2) = '0'   and
                (A1 or A1) = '1'   and
                (A1 or A2) = '1'   and
                (A2 or A1) = '1'   and
                (A2 or A2) = '0'   and
                (A1 xor A1) = '0'   and
                (A1 xor A2) = '1'   and
                (A2 xor A1) = '1'   and
                (A2 xor A2) = '0'   and
                (A1 nand A1) = '0'   and
                (A1 nand A2) = '1'   and
                (A2 nand A1) = '1'   and
                (A2 nand A2) = '1'   and
                (A1 nor A1) = '0'   and
                (A1 nor A2) = '0'   and
                (A2 nor A1) = '0'   and
                (A2 nor A2) = '1'   and
                (not A1) = '0'      and
                (not A2) = '1')
      report "***FAILED TEST: c07s02b01x00p02n02i01975 - BIT type truth table test failed." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c07s02b01x00p02n02i01975arch;
