library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

-- Documentation before pack_1
package pack_1 is
	-- Global constant const_1
	constant const_1 : boolean := false;

end package;

package body pack_1 is
	constant const_2 : boolean := true;

end package body;
