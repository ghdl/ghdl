package pkgb is
  constant b : natural := 2;
end;
