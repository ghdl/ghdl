package attrs_pkg is

  attribute ent_name: string;
  attribute ent_type: string;
  attribute ent_stat: integer;

  attribute arc_name: string;
  attribute arc_type: string;
  attribute arc_stat: integer;

end package;
