entity tb is
end entity;

architecture h of tb is
begin
  t:entity k't port map(0);
end architecture;
