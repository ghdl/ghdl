library ieee;use ieee.std_logic_1164;use ieee.numeric_std.all;entity hello is
port(c:std'l;t:d(0));end hello;architecture behav of h is
signal v:d(0);begin
process(c)begin
if(0)then
if 0='0'then
s;end if;end if;end process;end behav;