
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1478.vhd,v 1.2 2001-10-26 16:30:10 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c08s08b00x00p04n01i01478ent IS
END c08s08b00x00p04n01i01478ent;

ARCHITECTURE c08s08b00x00p04n01i01478arch OF c08s08b00x00p04n01i01478ent IS

BEGIN
  TESTING: PROCESS
    type i_array_type is array (1 to 5) of integer;
    variable a1 : i_array_type := (others => 0);
  BEGIN

    case a1 is                        -- illegal, must be discrete
      when 0 =>
        assert false
          report "Array allowed as case expression."
          severity note ;
      when others =>
        assert false
          report "Array allowed as case expression."
          severity note ;
    end case;

    assert FALSE 
      report "***FAILED TEST: c08s08b00x00p04n01i01478 - Array type is not allowed in expression." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c08s08b00x00p04n01i01478arch;
