architecture arch of ent is
  --  Comment for :b2:
  signal b2 : bit;
begin
end arch;
