entity e is
  generic(type t);
  signal w:integer range 0 to t(0);
end;
