entity attr is
end attr;

architecture behav of attr is
  attribute my_attr : ;
begin
end behav;
