package--
function is
if)h';