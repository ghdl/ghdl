architecture arch of ent is
  signal b1 : bit;

  --  Comment
  signal b2 : bit;
begin
end arch;
