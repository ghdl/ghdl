%%d%