library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package TestPkg is
  type ARecType is record
    A : unsigned(7 downto 0) ;
  end record ARecType ; 

end package TestPkg ; 
