
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1158.vhd,v 1.2 2001-10-26 16:30:03 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

package c06s06b00x00p02n01i01158pkg is
  type    I1    is range 1 to 5;
  subtype    I11    is I1 range 2 to 4;
  type    A1    is array (I1 range 2 to 4) of BOOLEAN;
end c06s06b00x00p02n01i01158pkg;

use work.c06s06b00x00p02n01i01158pkg.all;
ENTITY c06s06b00x00p02n01i01158ent IS
  generic (V_all : A1 := (true,false,true));
  port    (PT: BOOLEAN);
END c06s06b00x00p02n01i01158ent;

ARCHITECTURE c06s06b00x00p02n01i01158arch OF c06s06b00x00p02n01i01158ent IS

BEGIN
  TESTING: PROCESS
    variable  V      : boolean;
    attribute AT1    : A1;
    attribute AT1    of V : variable is V_all;
    variable  k    : integer := 0;
  BEGIN
    if I11'BASE'Left = 1 then
      k := 5;
    end if;
    assert NOT( k=5 )
      report "***PASSED TEST: c06s06b00x00p02n01i01158"
      severity NOTE;
    assert ( k=5 )
      report "***FAILED TEST: c06s06b00x00p02n01i01158 - The prefix of an attribute name may be a selected name." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c06s06b00x00p02n01i01158arch;
