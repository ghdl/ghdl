package pkg2 is
  generic (
    function func (a: integer) return natupac of integer
    );
end pkg2;
