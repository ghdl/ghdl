configuration cfg2 of e2 is
  -- comments in design units (python doc-string style)
  -- might be multi line
  for a2
  end for;
end configuration;
