package function is;X';