entity hello is
end hello;

architecture behav of hello is
begin
  << constant .h.x : bit >>;
end behav;
