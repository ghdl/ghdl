package p is
  function A return yy;
  function B return p'xx;
end;

