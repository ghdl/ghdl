
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc3016.vhd,v 1.2 2001-10-26 16:29:50 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

library WORK, STD;
use STD.STANDARD.all;   -- No_failure_here

ENTITY c11s02b00x00p05n02i03016ent IS
END c11s02b00x00p05n02i03016ent;

ARCHITECTURE c11s02b00x00p05n02i03016arch OF c11s02b00x00p05n02i03016ent IS
  signal BV : BIT_VECTOR(0 to 7);
BEGIN
  TESTING: PROCESS
  BEGIN
    BV <= "01010111" after 5 ns;
    wait for 10 ns;
    assert NOT( BV = "01010111" )
      report "***PASSED TEST: c11s02b00x00p05n02i03016"
      severity NOTE;
    assert ( BV = "01010111" )
      report "***FAILED TEST: c11s02b00x00p05n02i03016 - Library clause should appear as part of a context clause at the beginning of a design unit."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c11s02b00x00p05n02i03016arch;
