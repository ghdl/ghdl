
-- Copyright (C) 2002 Morgan Kaufmann Publishers, Inc

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

entity limiter is
  generic ( limit_high : real := 4.8;	 -- upper limit
            limit_low : real := -4.8 );  -- lower limit
  port ( quantity input : in real;
         quantity output : out real);					
end entity limiter;

----------------------------------------------------------------

architecture simple of limiter is
  constant slope : real := 1.0e-4;
begin

  if input > limit_high use    -- upper limit exceeded, so limit input signal
    output == limit_high + slope*(input - limit_high);
  elsif input < limit_low use  -- lower limit exceeded, so limit input signal
    output == limit_low + slope*(input - limit_low);
  else		               -- no limit exceeded, so pass input signal as is
    output == input;
  end use;

  break on input'above(limit_high), input'above(limit_low);

end architecture simple;
