package n is
  generic(package g is new w generic map(<>));
  function t return l;
end;
