
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc891.vhd,v 1.2 2001-10-26 16:30:01 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c10s02b00x00p02n02i00891ent IS
END c10s02b00x00p02n02i00891ent;

ARCHITECTURE c10s02b00x00p02n02i00891arch OF c10s02b00x00p02n02i00891ent IS
  type rec_typ is RECORD
                    -- immediate scope
                    r,g,b : real;
                  end record;
BEGIN
  TESTING: PROCESS
    -- extended scope
    variable electron_gun : rec_typ := ( 0.25, 0.5, 1.0 );
  BEGIN
    assert NOT(   electron_gun.r   = 0.25   and
                  electron_gun.g   = 0.5   and
                  electron_gun.b   = 1.0   ) 
      report "***PASSED TEST: c10s02b00x00p02n02i00891"
      severity NOTE;
    assert (   electron_gun.r   = 0.25   and
               electron_gun.g   = 0.5   and
               electron_gun.b   = 1.0   ) 
      report "***FAILED TEST: c10s02b00x00p02n02i00891 - The scope of the declaration that occurs immediately within a record type declaration extends beyond the immediate scope"
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c10s02b00x00p02n02i00891arch;
