
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2854.vhd,v 1.2 2001-10-26 16:29:49 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c13s10b00x00p03n01i02854ent IS
END c13s10b00x00p03n01i02854ent;

ARCHITECTURE c13s10b00x00p03n01i02854arch OF c13s10b00x00p03n01i02854ent IS
  constant   one    : integer := 16:E:E1;
  constant   two    : integer := 16#E#E1;
  constant   three   : integer := 16#FF#;
  constant   four   : integer := 16:FF:;
  constant   five   : integer := 2#1110_0000#;
  constant   six   : integer := 2:1110_0000:;
  constant   seven   : integer := 8#776#;
  constant   eight   : integer := 8:776:;
BEGIN
  TESTING: PROCESS
  BEGIN
    wait for 5 ns;
    assert NOT(    one=two    and 
                   three=four    and 
                   five=six    and 
                   seven=eight    )
      report "***PASSED TEST: c13s10b00x00p03n01i02854"
      severity NOTE;
    assert (    one=two    and 
                three=four    and 
                five=six    and 
                seven=eight    )
      report "***FAILED TEST: c13s10b00x00p03n01i02854 - Colon(:) can replace the sharp character(#) in based literal definition."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c13s10b00x00p03n01i02854arch;
