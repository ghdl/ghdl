library ieee;
use ieee.math_real.all;

entity test_64bit is

end entity test_64bit;

architecture sim of test_64bit is
begin

end architecture sim;
