library ieee;use ieee.numeric_std.all;use ieee.std_logic_1164.all;entity t is generic(e:boolean:=false);port(l:std'c);end;architecture a of g is type y is array(0)of t;signal m:n;begin
y<='0'when(0)else'0'when(0)and(0);process(l)begin
if(0)then if 0 then(0)<=0;end if;if 0 then if 0 then end if;end if;end if;end process;end;