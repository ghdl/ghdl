architecture arch of ent is
  --  Comment for :arch:
  --  Again for :arch:

  --  Also for :arch:

  --  But for :b1:
  signal b1 : bit;
begin
end arch;
