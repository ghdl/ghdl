library ieee;
use ieee.std_logic_1164.all;

entity badloc is
  constant v : std_logic_vector := b"01_X0";
end;
