entity repro6 is
end;

architecture behav of repro6 is
  type states_t is (s0, s1, s2);
  subtype st1 is states_t range s0 to s1;
begin
end behav;
