package p is
  type state_t is
    (
      s1,
      s2,
      --  Comment for :s3:
      s3);
end p;
