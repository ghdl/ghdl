architecture if''e';