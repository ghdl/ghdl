entity ent is
end ent;

architecture arch of ent is
begin
process begin report "Hello"; wait; end process;
end;
