library ieee ;
use ieee.std_logic_1164.all;

entity myentity is
end myentity;

architecture arch of myentity is
begin
end arch; 
