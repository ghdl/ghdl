package gen0 is
generic(v:natural:=0);function get return natural;end gen0;package body gen0 is
function get return natural is
begin
return+0;end get;end gen0;package gen0 is
generic(package p is new k'g generic map(<>));function t return l;end gen0;package n is use p;end;package g is new k;package p is new n generic map(0);entity b is
end;architecture behav of b is
begin a;end behav;