-- My comment �� îOD:x

entity ent is
end;
