entity inst1 is
end;

architecture behav of inst1 is
begin
   ins : entity ;
end behav;
