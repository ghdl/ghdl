context a is
  library ieee;
  context b is
  end;
end;
