library ieee;use ieee.numeric_std.all;use ieee.std_logic_1164.all;entity g is generic(type m;e:integer:=0;e0:boolean:=false);port(l:std'c);end;architecture a of g is type e;signal r:r range 0 to 0;signal r:r range 0 to 0;signal m:e;signal d:n;begin d(0);process(a)begin
if(0)then if 0 then m<=0;end if;if 0 then
elsif 0 then if 0 then r;end if;end if;end if;end process;end;