
-- Copyright (C) 2002 Morgan Kaufmann Publishers, Inc

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

library ieee_proposed;  use ieee_proposed.electrical_systems.all;
                        
entity quad_opamp is
  port ( terminal plus_in, minus_in, output : electrical_vector(1 to 4) );
end entity quad_opamp;

----------------------------------------------------------------

architecture slew_limited of quad_opamp is
  
  constant gain : real := 50.0;
  quantity v_in across plus_in to minus_in;
  quantity v_out across i_out through output;
  quantity v_amplified : real_vector(1 to 4);
        
begin

  v_amplified(1) == gain * v_in(1);
  v_amplified(2) == gain * v_in(2);
  v_amplified(3) == gain * v_in(3);
  v_amplified(4) == gain * v_in(4);
  
  real_vector(v_out) == v_amplified'slew(1.0e6,-1.0e6);
  
end architecture slew_limited;
