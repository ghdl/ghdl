
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc970.vhd,v 1.2 2001-10-26 16:30:29 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c06s03b00x00p05n01i00970ent IS
END c06s03b00x00p05n01i00970ent;

ARCHITECTURE c06s03b00x00p05n01i00970arch OF c06s03b00x00p05n01i00970ent IS

BEGIN
  TESTING: PROCESS
    type x is
      record
        y : integer;
        z : boolean;
      end record;
    type a is
      record
        b : real;
        c : integer;
      end record;
    variable r : a;
    variable p : x;
  BEGIN
    p.b := 1;   -- the prefix is not of an appropriate type as the 'p' does
    a.y := 1;   -- not have field 'b' and 'a' does not have field 'y'.   
    assert FALSE 
      report "***FAILED TEST: c06s03b00x00p05n01i00970 - Prefix is not apropraite for the type of the suffix." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c06s03b00x00p05n01i00970arch;
