-- comments before design units :cfg1:
-- might be multiline :cfg1:
configuration cfg1 of e1 is
  for a1
  end for;
end configuration;
