
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1210.vhd,v 1.2 2001-10-26 16:29:39 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c08s01b00x00p25n01i01210ent IS
END c08s01b00x00p25n01i01210ent;

ARCHITECTURE c08s01b00x00p25n01i01210arch OF c08s01b00x00p25n01i01210ent IS
  signal T1 : BIT := '0';
BEGIN
  TESTING: PROCESS
  BEGIN
    T1 <= '1' after 15 ns;
    wait on T1 until (T1 = '1');
    assert NOT( T1 = '1' )
      report "***PASSED TEST: c08s01b00x00p25n01i01210"
      severity NOTE;
    assert ( T1 = '1' )
      report "***FAILED TEST: c08s01b00x00p25n01i01210 - Process resumes execution when the condition clause in a wait statement is met"
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c08s01b00x00p25n01i01210arch;
