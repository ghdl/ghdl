package p is
  --  Comment for the record
  type rec is record
    a : bit;
    b : bit;
  end record;
end p;
