entity st2 is
end;

architecture arch of st2 is
  subtype mypos is natural range -1 to 5;
  subtype my2 is mypos range 2 to 3;
begin
end arch;
