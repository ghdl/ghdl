context ctx2 is
  -- comments in design units (python doc-string style)
    -- might be multi line
end context;

