entity top is
end top;
