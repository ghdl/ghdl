entity e is
end;

architecture a of e is
  constant a : real := 1000.0 / 100;
  constant b : time := 1000.0 / 100 * 10 ps;
begin
end;
