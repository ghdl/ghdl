entity begin restrict[*to 0