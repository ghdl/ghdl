
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1068.vhd,v 1.2 2001-10-26 16:30:06 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c06s04b00x00p03n04i01068ent IS
END c06s04b00x00p03n04i01068ent;

ARCHITECTURE c06s04b00x00p03n04i01068arch OF c06s04b00x00p03n04i01068ent IS

BEGIN
  TESTING: PROCESS
    variable str : string(1 to 20) := "This is string check";
  BEGIN
    if str(21) = 'T' then  -- illegal as 21 does not belong to the index
      -- range of str.
    end if;
    assert FALSE 
      report "***FAILED TEST: c06s04b00x00p03n04i01068 - Index value should belong to the range of the corresponding index range of the array." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c06s04b00x00p03n04i01068arch;
