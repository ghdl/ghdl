use work.a.all;

package b is
end package b;
