package--
function(0is;r';