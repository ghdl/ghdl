entity top is
end top;

use work.vc_fakeram_pkg;
architecture behav of top is
begin
end behav;
