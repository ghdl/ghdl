package function begin if t X';