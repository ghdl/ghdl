package t is
  type arr is array (natural range 0 to 7) of bit;
  subtype arridx is arr'range;
end t;
