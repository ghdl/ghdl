package p is
  --  Comment for :vec:
  type vec is array(natural) of bit_vector(0 to 1);
end p;
