entity package