package function begin n';