library ieee;
use ieee.std_logic_1164.all;

entity id2 is
  port (a_, b, ck : std_logic);
end;

architecture behav of id2 is
begin
end behav;
