package function begin--
X';