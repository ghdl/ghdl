library ieee;
use ieee.UPF.all;

entity test is
end entity;
