package arr_err1 is
  type t_slv32_x3 is array(1 tnatural range <>) of bit_vector(31 downto 0);
end arr_err1;

