package p is
  function log2(
    -- we also want to document parameters too
    param1 : integer;
    param2 : boolean
    ) return natural;
end p;


