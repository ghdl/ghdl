package repro is
  type array2d is array( integer range 0 to 7, integer range 14 downto 1)
  of natural;

  constant cst : array2d :=
  (
       (1,1,1,1,1,1,1,1,1,1,1,1,1,1),
       (2,3,5,9,17,33,65,129,257,513,1025,2049,4097,1),
       (3,5,9,17,33,65,129,257,513,1025,2049,4097,1,1),
       (4,7,13,25,49,97,193,385,769,1537,3073,6145,4097,1),
       (5,9,17,33,65,129,257,513,1025,2049,4097,1,1,1),
       (6,11,21,41,81,161,321,641,1281,2561,5121,2049,4097,1),
       (7,13,25,49,97,193,385,769,1537,3073,6145,4097,1,1),
       (8,15,29,57,113,225,449,897,1793,3585,7169,6145,4097,1)
   );

end repro;
