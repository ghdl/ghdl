entity t2 is
end entity;

architecture a of t2 is
  constant SimulationTime_c  : time    := 0.0 ps;
begin
end;

