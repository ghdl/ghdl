architecture arch of ent is
  signal b1 : bit;  --  Comment for :b1:
begin
end arch;
