package repro2 is
  type rec1 is record
    wr : bit;
    dat : bit_vector(7 downto 0);
  end record;
end repro2;
