entity module is
    generic(

    );
end entity;
