architecture behav of tb is
begin
  assert false report "Hello world" severity note;
end behav;
