library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity test4 is
end entity ;

architecture arch of test4 is

    constant x : signed(15 downto 0) := to_signed(0, 17);
begin
end architecture ;
