
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc347.vhd,v 1.2 2001-10-26 16:29:53 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s02b01x00p15n01i00347ent IS
END c03s02b01x00p15n01i00347ent;

ARCHITECTURE c03s02b01x00p15n01i00347arch OF c03s02b01x00p15n01i00347ent IS
  type MEM is array(5 downto 0) of BIT;  -- No_failure_here
  signal S1 : MEM := "000000";
BEGIN
  TESTING: PROCESS
  BEGIN
    assert NOT(S1(4 downto 3) = "00")
      report "***PASSED TEST: c03s02b01x00p15n01i00347"
      severity NOTE;
    assert (S1(4 downto 3) = "00")
      report "***FAILED TEST: c03s02b01x00p15n01i00347 - The direction of the discrete range is the same as the direction of the range."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s02b01x00p15n01i00347arch;
