entity top is
end top;

use work.test_pkg;
architecture behav of top is
begin
end behav;
