use work.types_pkg.all;

package const_pkg is
    constant c : generic_type := (others => 5);
end package;
