package pkg is
end package;

context ctx is
  library lib;
  use lib.pkg.all;
end context;
