library ieee;use ieee.std_logic_1164;entity t is
port(s:std'l);end entity;architecture a of t is
begin	i;end architecture;library i;entity b is
end entity;architecture h of b is
signal n:r(0);signal s:s(0);begin process	begin
end process;t(0);end architecture;