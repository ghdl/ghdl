
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1719.vhd,v 1.2 2001-10-26 16:29:43 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c09s02b00x00p16n02i01719ent IS
END c09s02b00x00p16n02i01719ent;

ARCHITECTURE c09s02b00x00p16n02i01719arch OF c09s02b00x00p16n02i01719ent IS
  SUBTYPE bit_4 is bit_vector ( 0 to 3);
  SUBTYPE bit_8 is bit_vector ( 0 to 7);

  SIGNAL  s  : bit_8 := B"0000_0000";
  SIGNAL  s4 : bit_4;
  SIGNAL  s5 : bit_4;
BEGIN

  -- trigger only one element.
  s (6) <= '1' after 10 ns;

  TESTING: PROCESS(s(0 to 3))
  BEGIN
    assert (NOW <= 0 fs ) 
      report "***FAILED TEST: c09s02b00x00p16n02i01719 - This process should be inactive."
      severity ERROR;
  END PROCESS TESTING;

  p2 : PROCESS (s(3 to 6))
  begin
    assert NOT((s(3 to 6) = B"0001") and (NOW = 10 ns))
      report "***PASSED TEST: c09s02b00x00p16n02i01719 - This test is passed only is the FAILED assertion did not appear."
      severity NOTE;
  end process p2;


END c09s02b00x00p16n02i01719arch;
