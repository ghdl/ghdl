entity ent is
end;

architecture structural of ent is
  constant stillOk    : integer := -2147483599;
  constant underflows : integer := -2147483600;
begin
end;
