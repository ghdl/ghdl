package g0 is
  package is
  end package;
end package;
