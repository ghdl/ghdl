architecture behav of tb is
begin
  assert work.pkg2.get2 = 5;
end behav;
