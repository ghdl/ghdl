entity repro3 is
end;

architecture behav of repro3 is
  component comp is
  end component comp;
  constant d : time := 1 comp;
begin
end behav;
