package function begin--
n';