package allnl is
  constant cr_eol : integer := 0;
  constant lf_eol : integer := 0;constant crlf_eol : integer := 0;
  constant lfcr_eol : integer := 0;
end allnl;
