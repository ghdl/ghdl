
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2982.vhd,v 1.2 2001-10-26 16:29:50 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

package c02s05b00x00p01n01i02982pkg is
  type       tristate    is ('0','1','Z');
  subtype    bi       is integer range 1 to 2;
  constant    lowstate   : tristate:='0';
end c02s05b00x00p01n01i02982pkg;


ENTITY c02s05b00x00p01n01i02982ent IS
END c02s05b00x00p01n01i02982ent;

ARCHITECTURE c02s05b00x00p01n01i02982arch OF c02s05b00x00p01n01i02982ent IS
  use work.c02s05b00x00p01n01i02982pkg.all;
BEGIN
  TESTING: PROCESS
    variable locz:tristate   :='Z';
    variable loch:bi   :=2;
  BEGIN
    locz:=lowstate;
    loch:=1;
    wait for 5 ns;
    assert NOT( locz='0' and loch<2 )
      report "***PASSED TEST: c02s05b00x00p01n01i02982"
      severity NOTE;
    assert ( locz='0' and loch<2 )
      report "***FAILED TEST: c02s05b00x00p01n01i02982 - Package declaration syntax test failed."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c02s05b00x00p01n01i02982arch;
