entity tb is
end tb;
