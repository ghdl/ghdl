package p is
  --  Comment
  type vec is array(natural range <>) of bit_vector(0 to 1);
end p;
