package p2 is
  -- comments in design units (python doc-string style) :fail:
end package;
