library ieee;
use ieee.std_logic_1164.all;

package mixer_pkg is
    type sample_array is array (natural range <>) of std_logic_vector;
end package mixer_pkg;
