--  comment for :a2:
architecture a2 of e2 is
  -- comments in design units (python doc-string style) :a2:
  --:a2: might be multi line

  --  comment for :s:
  signal s : bit;
begin

end architecture;
