package nullrng is

  type my_empty_range is range -(-8) to 7;
  type my_small_range is range -8 to 7;

end;
