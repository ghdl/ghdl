entity t is
end;

architecture behav of t is
begin
  assert (1 + 1) * 1 = 2;
end behav;
