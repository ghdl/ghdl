package pkg is
  constant time_image : time'image(now);
end package;
