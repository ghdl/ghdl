entity test is end entity; 

architecture arch of test is 
  signal b:bit; 
  alias bit_base is bit'base; 
  -- alias b_stable is b'stable; 
begin 
end architecture; 
