entity hello is
end hello;

use work.pkg.all;
architecture behav of hello is
begin
  say_hello;
end behav;
