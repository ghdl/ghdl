library ieee;
use ieee.numeric_bit.all;

entity t2 is
end;

architecture behav of t2 is
begin
  assert rising_edge('1');
end behav;
