library ieee;
use ieee.std_logic_1164.all;
entity test is
    port (
        clk     : in  std_logic
    );
end entity test;
architecture rtl of test is
begin
end architecture rtl;
