entity tb1 is
end tb1;

use work.pkg1.all;

architecture behav of tb1 is
begin
end behav;
