-- Author:  Patrick Lehmann
-- License: MIT
--
-- undocumented
--
context StopWatch_ctx is
	library lib_Utilities;
	context lib_Utilities.Utilities_ctx;

	library lib_Display;
	use     lib_Display.Display_pkg.all;

	use work.StopWatch_pkg.all;
end context;
