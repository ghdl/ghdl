entity st1 is
end;

architecture arch of st1 is
  subtype mypos is natural range -1 to 5;
begin
end arch;
