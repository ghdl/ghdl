entity hello is
end hello;
