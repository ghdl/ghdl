package pkg is
end pkg;
