package aa is
constant a : integer_vector(0 to 1) := (0, 1);
constant b : integer_vector(0 to 0) := a(integer range 0 to 0);
end package aa;
