CONTEXT is
context is