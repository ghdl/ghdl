entity t1 is
end entity;

architecture a of t1 is
  constant SimulationTime_c  : time    := 0 fs;
begin
end;

