entity nochoice is
end;

architecture behav of nochoice is
  constant n : natural := 5;
begin
  process
  begin
    case n is
    end case;
  end process;
end behav;
