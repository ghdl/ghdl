-- comments before design units (javadoc / .net documentation style)
-- might be multiline
entity e1 is
end entity;

-- comments before design units
-- might be multiline
architecture a1 of e1 is
begin
end architecture;

-- comments before design units
-- might be multiline
package p1 is
end package;

-- package body should be supported too to keep parity, but I have currently no usecase for it.

-- comments before design units
-- might be multiline
context ctx1 is
end context;

-- comments before design units
-- might be multiline
configuration cfg1 of e1 is
  for a1
  end for;
end configuration;


library ieee;
use ieee.std_logic_1164.all;

entity e2 is
  -- comments in design units (python doc-string style)
    -- might be multi line
    generic (
      -- comment before a generic
        -- might be multiline
        constant FREQUENCY : positive;
      constant BITS      : positive; -- comment after a generic are mostly single line,
                                       -- but could be multi line too
        -- in case comment is before and after
        constant DEBUG     : boolean   -- the after has presidence
    );
    port (
      signal Clock : in std_logic    -- same as for generics
    );
end entity;

architecture a2 of e2 is
  -- comments in design units (python doc-string style)
    -- might be multi line
begin

end architecture;

-- As packages define public elements like constants, types and sub-programs, we are intrested in such documentation too.
package p2 is
  -- comments in design units (python doc-string style)
    -- might be multi line

    -- comment before
    constant DEBUG : boolean := TRUE;
    constant SYNC_STAGES : positive := 3; -- comment after

    -- comment before
    type AType1 is array(natural range <>) of bit;
    type AType2 is array(natural range <>) of bit; -- comment after

    -- same applies to subtype, alias, attributes, ...

    -- comment before
    type RType is record
        -- xor comment inside

        -- per element comment before (note the comment "block" is separated by newlines)
        elem1 : integer;
        elem2 : integer; -- per element comment behind
    end record;

    -- as functions are longer in definitions, it might be written before
    function log2(param : positive) return natural;

    function log2(
        -- otoh, we also want to document parameters too (similar to a record with comments)

      -- comment before
      param1 : integer;
        param2 : boolean  -- comment after
    ) return natural;

    -- this applies to procedures as well.



end package;

context ctx2 is
  -- comments in design units (python doc-string style)
    -- might be multi line
end context;

configuration cfg2 of e2 is
  -- comments in design units (python doc-string style)
  -- might be multi line
  for a2
  end for;
end configuration;







-- This should allow for any kind of documentation style and embedded documentation language.
-- A real implementation might use similar rules are Python+docutils+Sphinx. Here we would e.g.
-- document a function either before (or inside) a function declaration and use the
--   :arg name: description
-- syntax.


-- Package `math` provides math extensions not provided by the IEEE packages.
package math is
    -- Computes the logarith to base 2.
    --
    -- :arg param: Input value
    -- :returns:   Logarithm
    function log2(param : positive) return natural;
end package;
