-- comments before design units :a1:
-- might be multiline :a1:
architecture a1 of e1 is
begin
end architecture;
