package n is
  function t return n;
end;
package body n is
  function get return l is
  begin
  end get;
end;

package n is
  generic(package g is new w generic map(<>));
  function t return l;
end;

package body gen0 is
  use p;
  function g return l is
  begin
  end;
end gen0;

package b is
end;

architecture beha0 of b is
begin
end beha0;
