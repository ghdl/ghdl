architecture restrict[*9000000000