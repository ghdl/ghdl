library ieee;
use ieee.std_logic_1164.all;

package repro is
  alias reg_Acc : std_logic_vector(3 downto 0) is "0111";
end repro;
