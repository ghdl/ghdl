library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package compa_pkg is

type test_rec is record
	a	: std_logic_vector;
	b	: std_logic_vector;
end record;


end package;
