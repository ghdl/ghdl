library ieee;
use ieee.std_logic_1164.all;

entity quote1 is
  constant v : std_logic_vector := b%0_10";
end;
