
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc112.vhd,v 1.2 2001-10-26 16:30:06 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c04s03b02x00p29n06i00112ent IS
  port (   S1 : out BIT_VECTOR(0 to 3) := "1011";
           S2 : out BIT := '1') ;
END c04s03b02x00p29n06i00112ent;

ARCHITECTURE c04s03b02x00p29n06i00112arch OF c04s03b02x00p29n06i00112ent IS
  signal S3 : BIT;
BEGIN

  S3    <= S2 after 20 ns;      --Failure here

  TESTING: PROCESS
  BEGIN
    assert FALSE
      report "***FAILED TEST: c04s03b02x00p29n06i00112 - Interface object of mode out cannot be read."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c04s03b02x00p29n06i00112arch;
