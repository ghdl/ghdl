entity str is
end str;

architecture behav of str is
begin
  process
  begin
    null;
    "abc";
    null;
  end process;
end behav;
