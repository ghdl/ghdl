entity reserved1 is
end reserved1;

architecture behav of reserved1 is
  signal quantity : bit;
begin
  process
  begin
    wait;
  end process;
end behav;
