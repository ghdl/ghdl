
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc943.vhd,v 1.2 2001-10-26 16:30:02 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c06s01b00x00p08n01i00943ent IS
END c06s01b00x00p08n01i00943ent;

ARCHITECTURE c06s01b00x00p08n01i00943arch OF c06s01b00x00p08n01i00943ent IS

BEGIN
  TESTING: PROCESS
    variable V1 : BIT_VECTOR(0 to 5);     -- No_failure_here
  BEGIN
    assert NOT( V1="000000" )
      report "***PASSED TEST: c06s01b00x00p08n01i00943"
      severity NOTE;
    assert ( V1="000000" )
      report "***FAILED TEST: c06s01b00x00p08n01i00943 - The name must be a simple name, an operator symbol, a selected name, an indexed name, a slice name, or an attribute name."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c06s01b00x00p08n01i00943arch;
