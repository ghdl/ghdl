
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc3104.vhd,v 1.2 2001-10-26 16:30:25 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c05s01b00x00p16n02i03104ent IS
  port    (PT:BOOLEAN);
  attribute AT1 : integer;
  attribute AT1 of ch0501_P01602_02_ent : entity is 1.2;  --  Failure_here
  --ERROR:  Specification expression is not the same type as attribute declaration
END c05s01b00x00p16n02i03104ent;

ARCHITECTURE c05s01b00x00p16n02i03104arch OF c05s01b00x00p16n02i03104ent IS

BEGIN
  TESTING: PROCESS
  BEGIN
    assert FALSE
      report "***FAILED TEST: c05s01b00x00p16n02i03104 - Specification expression is not of the same type as attribute specification."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c05s01b00x00p16n02i03104arch;
