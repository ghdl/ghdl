
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2565.vhd,v 1.2 2001-10-26 16:29:48 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c07s04b01x00p08n01i02565ent IS
END c07s04b01x00p08n01i02565ent;

ARCHITECTURE c07s04b01x00p08n01i02565arch OF c07s04b01x00p08n01i02565ent IS
  SUBTYPE s10 IS STRING (1 TO 4);

  ATTRIBUTE attr1 : INTEGER;
--
  ATTRIBUTE attr1 OF s10 : SUBTYPE IS 4;
BEGIN
  TESTING: PROCESS
    VARIABLE v : s10;
  BEGIN
--
--      The expressions in a named assocition list of more than 1 element
--      must be locally static.
--
    v := (1 | s10'attr1 => 'a', OTHERS => 'b' );
    wait for 5 ns;
    assert NOT( v="abba" )
      report "***PASSED TEST: c07s04b01x00p08n01i02565"
      severity NOTE;
    assert ( v="abba" )
      report "***FAILED TEST: c07s04b01x00p08n01i02565 - Bad value for named aggregate."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c07s04b01x00p08n01i02565arch;
