library ieee ;
use ieee.std_logic_1164.all;

entity myentity is
  port (
    inout1: inout std_logic_vector(9 downto 1) := "10ZWLH-UX"
    );
end myentity;

architecture arch of myentity is
begin
end arch;
