library IEEE;use IEEE.numeric_std.all;entity tb is
end;architecture behavioral of tb is
subtype int01 is integer range-0**(-1)to(0);type a is array(0)of i;function A(v:l)return r is variable p:d(0);begin e(0)(0);r((0));end;begin
process
variable t:t;variable tmp:int01;begin	tmp:=0;end process;end behavioral;