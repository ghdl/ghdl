package p is
  type rec is record
    a : bit; --  Comment for :a:
    --  Also for :a:
    b : bit;
  end record;
end p;
