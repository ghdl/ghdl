entity repro2 is
end;

architecture behav of repro2 is
  constant c : string := "hello";
  constant d : time := 1.5e2 c'length;
begin
end behav;
