package body function begin 0package