package pkg1 is new work.gen1;
