
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc911.vhd,v 1.2 2001-10-26 16:30:02 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

entity c10s03b00x00p07n01i00911ent_a is
end c10s03b00x00p07n01i00911ent_a;

architecture c10s03b00x00p07n01i00911arch_a of c10s03b00x00p07n01i00911ent_a is
begin
  TESTING : PROCESS
  BEGIN
    assert FALSE 
      report "***PASSED TEST: c10s03b00x00p07n01i00911"
      severity NOTE;
    wait;
  END PROCESS TESTING;
end c10s03b00x00p07n01i00911arch_a;


ENTITY c10s03b00x00p07n01i00911ent IS
END c10s03b00x00p07n01i00911ent;

ARCHITECTURE c10s03b00x00p07n01i00911arch OF c10s03b00x00p07n01i00911ent IS
  component device
  end component;

  -- selected use of configuration primary unit
  for all : device use entity work.c10s03b00x00p07n01i00911ent_a(c10s03b00x00p07n01i00911arch_a);
BEGIN
  instance : device;
END c10s03b00x00p07n01i00911arch;
