
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc272.vhd,v 1.2 2001-10-26 16:29:49 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s01b03x00p06n01i00272ent IS
END c03s01b03x00p06n01i00272ent;

ARCHITECTURE c03s01b03x00p06n01i00272arch OF c03s01b03x00p06n01i00272ent IS
  type small is range 0 to 2_000_000_000      --   < 2**31-1
    units
      lu;
    end units;
BEGIN
  TESTING: PROCESS
    variable   smaller : small;
  BEGIN
    smaller := 2000000000 lu;
    wait for 5 ns;
    assert NOT( smaller = 2000000000 lu ) 
      report "***PASSED TEST: c03s01b03x00p06n01i00272" 
      severity NOTE;
    assert ( smaller = 2000000000 lu ) 
      report "***FAILED TEST: c03s01b03x00p06n01i00272 - Large physical type declaration test failed."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s01b03x00p06n01i00272arch;
