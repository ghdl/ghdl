package body gen2 is
  use pkg.all;
  
  function get2 return natural is
  begin
    return get;
  end get2;
end gen2;
