library ieee;
use ieee.std_logic_signed;

entity tb is
end tb;
