entity reserved4 is
end;

architecture behav of reserved4 is
  signal xnor : bit;
begin
  process
  begin
    wait;
  end process;
end behav;
