package types_pkg is
    type t_symbol is (NARROW_SYMBOL, REGULAR_SYMBOL, WIDE_SYMBOL);
end package;
