package pkg1 is
  constant c : natural := 12;
end;
