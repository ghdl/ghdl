
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1146.vhd,v 1.2 2001-10-26 16:30:06 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c06s05b00x00p05n02i01146ent IS
END c06s05b00x00p05n02i01146ent;

ARCHITECTURE c06s05b00x00p05n02i01146arch OF c06s05b00x00p05n02i01146ent IS

BEGIN
  TESTING: PROCESS
    TYPE A IS ARRAY (NATURAL RANGE <>) OF INTEGER;
    SUBTYPE A6 IS A (1 TO 6);
    SUBTYPE A8 IS A (1 TO 8);
    FUNCTION func1 RETURN A6 IS
    BEGIN
      RETURN (1,2,3,4,5,6);
    END;
    VARIABLE ReturnValue : A8;
  BEGIN
    ReturnValue := func1(1 TO 8);
    assert FALSE 
      report "***FAILED TEST: c06s05b00x00p05n02i01146 - The bounds of the discrete range does not belong to the index range of the prefixing array." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c06s05b00x00p05n02i01146arch;
