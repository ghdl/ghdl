entity crash_Tb is
end;

use work.crash_pkg.all;
architecture behav of crash_tb is
begin
end behav;
