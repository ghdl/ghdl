package gen1 is
  generic (v : natural := 5);

  function get return natural;
end gen1;
