package pkg3 is
  function f (a : integer) return integer;
  function f (a : integer) return integer is
  begin
   return 1;
  end f;
end pkg3;
