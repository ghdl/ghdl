package p is

  constant c : natural := 1;

  --  Comment for :rec:
  type rec is record
    a : bit;
    b : bit;
  end record;
end p;
