library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

vunit const_test_vunit (const_test(rtl))
{
    constant depth : positive := 2**addr_width;
}
