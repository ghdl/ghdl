entity hello is
  port(c:s't bit_vector(0));
end hello;
