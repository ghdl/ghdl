
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1797.vhd,v 1.2 2001-10-26 16:30:12 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c07s01b00x00p02n01i01797ent IS
END c07s01b00x00p02n01i01797ent;

ARCHITECTURE c07s01b00x00p02n01i01797arch OF c07s01b00x00p02n01i01797ent IS
  -- architecture declaration section
BEGIN
  -- architecture statement part
  TESTING: PROCESS
  BEGIN
    -- testcase code
    Assert FALSE
      Report "***PASSED TEST: c07s01b00x00p02n01i01797"
      Severity NOTE;
    -- testcase code
    Assert FALSE
      Report "***FAILED TEST: c07s01b00x00p02n01i01797"
      Severity ERROR;
    wait; -- forever
  END PROCESS TESTING;
END c07s01b00x00p02n01i01797arch;

-- CONFIGURATION c07s01b00x00p02n01i01797cfg OF c07s01b00x00p02n01i01797ent IS
--     FOR c07s01b00x00p02n01i01797arch
--     END FOR;
-- END c07s01b00x00p02n01i01797cfg;

