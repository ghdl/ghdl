package function is;i';