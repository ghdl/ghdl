library ieee;
use ieee.std_logic_1164.all;

entity e is
    generic (file f : integer);
end entity;

architecture a of e is
begin
end architecture;
