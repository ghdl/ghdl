package--
function is;n';