entity e is end entity;
architecture a of e is
  constant s1 :string := foreign'path;
  constant s2 :string := foreign'foreign;
begin
end architecture;
