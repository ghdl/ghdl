
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1643.vhd,v 1.2 2001-10-26 16:29:42 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

package c08s12b00x00p08n01i01643pkg is


  -- function declarations.
  function funcI  return INTEGER;
  function funcI2 return INTEGER;

end c08s12b00x00p08n01i01643pkg;

package body c08s12b00x00p08n01i01643pkg is

  function funcI return INTEGER is
  begin
    return ( 3 );
  end;

  function funcI2 return INTEGER is
  begin
    return ( 3  );
  end;

end c08s12b00x00p08n01i01643pkg;

use work.c08s12b00x00p08n01i01643pkg.all;
ENTITY c08s12b00x00p08n01i01643ent IS
END c08s12b00x00p08n01i01643ent;

ARCHITECTURE c08s12b00x00p08n01i01643arch OF c08s12b00x00p08n01i01643ent IS

BEGIN
  TESTING: PROCESS
  BEGIN
    assert NOT( funcI = 3 and funcI2 = 3)         
      report "***PASSED TEST: c08s12b00x00p08n01i01643"
      severity NOTE;
    assert ( funcI = 3 and funcI2 = 3)         
      report "***FAILED TEST: c08s12b00x00p08n01i01643 - "
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c08s12b00x00p08n01i01643arch;
