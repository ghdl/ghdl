package pkg is
 type e is (identifier, i2);
-- procedure identifier;
-- alias identifier_alias_fun is identifier[return integer];
 alias identifier_alias_proc is identifier[];
end package;
