library ieee;
use ieee.std_logic_1164.all;

entity bug2 is
end;

architecture behavior of bug2 is
begin
    std_logic(1 downto 0);
end behavior;
