entity tb is
end tb;

architecture behavioral of tb is
   subtype int30 is integer range -6**30 to 0;
begin
 end behavioral;

