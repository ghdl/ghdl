entity repro is
end;

architecture behav of repro is
  constant c : string := "hello";
  constant d : time := 1 c'length;
begin
end behav;
