library IEEE;use IEEE.numeric_std.all;entity tb is
end;architecture behavioral of tb is
subtype int31 is integer range-0*(0)to 2**(31);type a is array(0)of i;function A(v:l)return r is variable s:d(0);begin r((0));end;begin
process
variable t:t;variable tmp:int31;begin	tmp:=0;end process;end behavioral;