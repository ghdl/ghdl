
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2919.vhd,v 1.2 2001-10-26 16:30:24 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c02s01b01x02p06n01i02919ent IS
END c02s01b01x02p06n01i02919ent;

ARCHITECTURE c02s01b01x02p06n01i02919arch OF c02s01b01x02p06n01i02919ent IS
  procedure proc1 (signal x1 : bit; z1 : boolean);
  procedure proc1 (signal x1 : bit; z1 : boolean) is
  begin
    null;
  end proc1;
  signal b: bit_vector (4 downto 1);
BEGIN
  TESTING: PROCESS
    variable i : integer := 1;
  BEGIN
    proc1 (b(i), true);  -- Failure_here
    -- b(i) is not a static name.
    assert FALSE
      report "***FAILED TEST: c02s01b01x02p06n01i02919 - The actual signal associated with a signal parameter must be denoted by a static name."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c02s01b01x02p06n01i02919arch;
