package
function begin if a s';