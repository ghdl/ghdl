
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2200.vhd,v 1.2 2001-10-26 16:29:46 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c07s02b06x00p01n01i02200ent IS
END c07s02b06x00p01n01i02200ent;

ARCHITECTURE c07s02b06x00p01n01i02200arch OF c07s02b06x00p01n01i02200ent IS

BEGIN
  TESTING: PROCESS
    variable z : real := -0.01 / (1.0); -- z should be -0.01
  BEGIN
    assert NOT(z=-0.01)
      report "***PASSED TEST: c07s02b06x00p01n01i02200"
      severity NOTE;
    assert ( z=-0.01 )
      report "***FAILED TEST: c07s02b06x00p01n01i02200 - The  operators * and / are predefined for any integer type and any floating point type and have their convertional meaning."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c07s02b06x00p01n01i02200arch;
