package types_pkg is
    type generic_type is array(0 to 3) of integer;
end package;
