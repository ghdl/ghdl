d%