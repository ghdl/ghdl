`entity fum is
`end entity;
`
`architecture bul of fum is
`    begin
`    end architecture;
```
