entity ams1 is
end;

architecture behav of ams1 is
  nature electrical is real across real through ground reference;
  --  terminal nx : electrical;
  --  quantity energy : real;
begin
  process
  begin
    wait;
  end process;
end behav;
