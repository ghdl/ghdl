
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc511.vhd,v 1.2 2001-10-26 16:30:26 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s02b02x00p06n03i00511ent IS
END c03s02b02x00p06n03i00511ent;

ARCHITECTURE c03s02b02x00p06n03i00511arch OF c03s02b02x00p06n03i00511ent IS
  type R1 is record
               RE1: I1;
               RE2: RE1;  -- Failure_here
               -- ERROR - SEMANTIC ERROR: NAME OF RECORD ELEMENT CANNOT BE USED
               -- WITHIN THE RECORD TYPE DEFINITION
             end record;
BEGIN
  TESTING: PROCESS
  BEGIN
    assert FALSE 
      report "***FAILED TEST: c03s02b02x00p06n03i00511 - Name of record element cannot be used in the record type definition." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s02b02x00p06n03i00511arch;
