package p is

  constant c : natural := 1;

  --  Comment for the decl.
  constant c1 : natural := 3;
end p;
