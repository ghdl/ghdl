entity tab1 is
  port (
    p__1 : bit;
    abcd__2 : bit;
    bad_ : bit;
	ontab_ : bit;
        notab_ : bit;
    _err : bit;
    num : integer := 1_2_);
end tab1;
