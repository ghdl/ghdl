
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1705.vhd,v 1.2 2001-10-26 16:29:43 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c09s02b00x00p07n01i01705ent IS
END c09s02b00x00p07n01i01705ent;

ARCHITECTURE c09s02b00x00p07n01i01705arch OF c09s02b00x00p07n01i01705ent IS
  signal   S1 :    Bit;
  signal   S2 :    Bit;
BEGIN
  TESTING: PROCESS( S1 )
  BEGIN
    S1   <=   '1' after 10 ns;
  END PROCESS TESTING;

  TESTING1: PROCESS
  BEGIN
    S2   <=   '1' after 10 ns;
    wait on S2;
    assert NOT(S1=S2) 
      report "***PASSED TEST: c09s02b00x00p07n01i01705"
      severity NOTE;
    assert (S1=S2) 
      report "***FAILED TEST: c09s02b00x00p07n01i01705 - The process statement is assumed to contain an implicit wait statement if a sensitivity list appears following the reserved word process."
      severity ERROR;
    wait;
  END PROCESS TESTING1;

END c09s02b00x00p07n01i01705arch;
