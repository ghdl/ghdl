LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY json_format IS
END ENTITY json_format;

ARCHITECTURE rtl OF json_format IS
    SIGNAL clk : std_logic := '0';
BEGIN
    clk <= '1';

    main : PROCESS
    BEGIN
        WAIT;
    END PROCESS;

END ARCHITECTURE;
