-- Author:  Patrick Lehmann
-- License: MIT
--
-- A generic counter module used in the StopWatch example.
--
context StopWatch_ctx is
	library IEEE;
	use     IEEE.std_logic_1164.all,
	        IEEE.numeric_std.all;

	use work.StopWatch_pkg.all;
end context;
