
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc3022.vhd,v 1.2 2001-10-26 16:29:50 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

package c11s03b00x00p04n02i03022pkg is
  type T is (one,two,three,four);
  subtype SIN is INTEGER;
end c11s03b00x00p04n02i03022pkg;

use work.c11s03b00x00p04n02i03022pkg.all;
ENTITY c11s03b00x00p04n02i03022ent IS
END c11s03b00x00p04n02i03022ent;

ARCHITECTURE c11s03b00x00p04n02i03022arch OF c11s03b00x00p04n02i03022ent IS
  signal S1 : T;      -- type T should be visible
  signal S2 : SIN;    -- subtype SIN should be visible
  signal S3 : REAL;
BEGIN
  TESTING: PROCESS
  BEGIN
    S1 <= one;      --literal "one" should be visible
    S2 <= 1234;
    wait for 5 ns;
    assert NOT( S1 = one and S2 = 1234 )
      report "***PASSED TEST: c11s03b00x00p04n02i03022"
      severity NOTE;
    assert ( S1 = one and S2 = 1234 )
      report "***FAILED TEST: c11s03b00x00p04n02i03022 - A use clause should make certain declarations directly visible within the design unit."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c11s03b00x00p04n02i03022arch;
