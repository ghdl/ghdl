package bug_pkg is
  type t_zero_one is (zero, one);
end package bug_pkg;
