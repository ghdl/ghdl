
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc780.vhd,v 1.2 2001-10-26 16:30:27 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c01s01b01x02p11n01i00780ent IS
  port ( S : buffer bit );
END c01s01b01x02p11n01i00780ent;

ARCHITECTURE c01s01b01x02p11n01i00780arch OF c01s01b01x02p11n01i00780ent IS

BEGIN
  TEST : PROCESS
  BEGIN
    S <= bit'('1');
    wait for 15 ns;
  END PROCESS TEST;

  TESTING: PROCESS
  BEGIN
    S <= bit'('0'); -- Failure_here
    -- signal S of mode buffer is being
    -- driven by two sources one in each
    -- process. Signal S can be driven by
    -- only one source.
    -- This error will be indicated at elaboration time
    wait for 11 ns;
    assert FALSE
      report "***FAILED TEST: c01s01b01x02p11n01i00780 - A buffer port can have at most one source."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c01s01b01x02p11n01i00780arch;
