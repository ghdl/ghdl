
-- Copyright (C) 1996 Morgan Kaufmann Publishers, Inc

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: ap_a_ap_a_05.vhd,v 1.1.1.1 2001-08-22 18:20:47 paw Exp $
-- $Revision: 1.1.1.1 $
--
-- ---------------------------------------------------------------------

entity ap_a_05 is

end entity ap_a_05;


library ieee;  use ieee.std_logic_1164.all;

architecture test of ap_a_05 is

  signal a, b, y, x : std_ulogic;

begin

  -- code from book

  y <= a when x = '1' else
       b;

  -- end code from book

  x <= '0', '1' after 20 ns;
  a <= '0', '1' after 10 ns, '0' after 20 ns, '1' after 30 ns;
  b <= '0', '1' after 15 ns, '0' after 25 ns, '1' after 35 ns;

end architecture test;

