
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc779.vhd,v 1.2 2001-10-26 16:30:27 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c01s01b01x02p11n02i00779ent_a IS
  port (c2 : buffer Bit);
END c01s01b01x02p11n02i00779ent_a;

ARCHITECTURE c01s01b01x02p11n02i00779arch_a OF c01s01b01x02p11n02i00779ent_a IS
BEGIN
END c01s01b01x02p11n02i00779arch_a;



ENTITY c01s01b01x02p11n02i00779ent IS
  port(P2 : buffer Bit);
END c01s01b01x02p11n02i00779ent;

ARCHITECTURE c01s01b01x02p11n02i00779arch OF c01s01b01x02p11n02i00779ent IS
  component c01s01b01x02p11n02i00779ent_b
    port (C2 : buffer Bit);
  end component;
  for L : c01s01b01x02p11n02i00779ent_b use entity work.c01s01b01x02p11n02i00779ent(c01s01b01x02p11n02i00779arch) port map (C2);
BEGIN

  L : c01s01b01x02p11n02i00779ent_b port map (C2 => P2);

  TEST : Process
  begin
    P2 <= bit'('1');
    wait for 15 ns;
  end process TEST;

  TESTING: PROCESS
  BEGIN
    P2 <= bit'('0');   -- Failure_here
    -- This error will be indicated at elaboration time.
    wait for 11 ns;
    assert FALSE
      report "***FAILED TEST: c01s01b01x02p11n02i00779 - Actual can have at most one source."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c01s01b01x02p11n02i00779arch;
