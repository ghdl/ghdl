
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc69.vhd,v 1.2 2001-10-26 16:29:59 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c04s03b01x02p07n05i00069ent IS
END c04s03b01x02p07n05i00069ent;

ARCHITECTURE c04s03b01x02p07n05i00069arch OF c04s03b01x02p07n05i00069ent IS
  signal S1 : BIT_VECTOR(0 to 3) := ("0101" and "0101");
BEGIN
  TESTING: PROCESS
  BEGIN
    wait for 10 ns;
    assert NOT(    S1(0)   = '0'   and
                   S1(1)   = '1'   and
                   S1(2)   = '0'   and
                   S1(3)   = '1'   )
      report "***PASSED TEST: c04s03b01x02p07n05i00069"
      severity NOTE;
    assert (    S1(0)   = '0'   and
                S1(1)   = '1'   and
                S1(2)   = '0'   and
                S1(3)   = '1'   )
      report "***FAILED TEST: c04s03b01x02p07n05i00069 - Each subelement of the value of the composite subtype is the default value of the corresponding subelement of the signal."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c04s03b01x02p07n05i00069arch;
