library ieee;
use ieee.std_logic_1164.all.common.workall;
entity icache is end;
