-- Author:  Patrick Lehmann
-- License: MIT
--
-- undocumented
--
context Display_ctx is
	library lib_Utilities;
	context lib_Utilities.Utilities_ctx;

	use work.Display_pkg.all;
end context;
