entity e is end entity;
architecture a of e is
 signal s :boolean;
begin
 assert not s;
end architecture;
