library ieee;
use ieee.std_logic_arith.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;

entity a is
end entity a;

architecture RTL of a is
begin
end architecture RTL;
