package p is
  type rec is record
    --  Comment for the first element.
    a : bit;
    b : bit;
  end record;
end p;
