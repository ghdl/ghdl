package p is
end p;
