�   a00 i0000000000 i0 a0000  000000 r0000 <>0l000��xi000;
use i00000000 i000;use i000.Sll;
u::::::::::::0s0 i000.s0d�o000000000000 y i000;
use 000.w00   0s�d  000���00000) packageb0;00:0s00_]  c;

00 c�t : ou000n00(0�w000 0)0B
et�.all;�
entityh0000�0 s000 o0 h000_ is
 s0000  �0:u0000000(0 downto 0);begin
   if r0
use 000.w00   )s�dsssssssssssssssspackage pkg0 is
� type s array (n000000 range <>, block, c0000_000000)
	v00000) packageb0;
e�d pkg0;use g000.pkg0.all;

package pkg0 is�  function fncal�
end k00nctio�  �n
  f00