library ieee;
use ieee.std_logic_1164.all;

entity e is
    port (i : in std_logic_vector(2 downto 0) := ('1','0'));
end entity;

architecture a of e is
begin
end architecture;
