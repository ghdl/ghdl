entity tb is
end;

use work.model_pkg.all;

architecture behav of tb is
begin
end;
