package p is

  constant c : natural := 1;

  --  Comment for the record
  type rec is record
    a : bit;
    b : bit;
  end record;
end p;
