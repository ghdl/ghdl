use work.p1.all;

package p1 is
  constant c : natural := 5;
end p1;
