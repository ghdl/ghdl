-- This is iso 8859-1 (latin-1) encoding. �l�ve.
-- Last chars of the last line are (hexa): e9 6c e8 76 65 2e

package p1 is
end p1;

