package p is

  constant c : natural := 1;

  --  Comment for the decl :c1:
  constant c1 : natural := 3;
end p;
