-- :e1: comments before design units (javadoc / .net documentation style)
-- :e1: might be multiline
entity e1 is
end entity;

-- :a1: comments before design units
-- :a1: might be multiline
architecture a1 of e1 is
begin
end architecture;
