package function begin--
�';