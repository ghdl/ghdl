
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2435.vhd,v 1.2 2001-10-26 16:29:47 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c07s03b02x02p01n02i02435ent IS
END c07s03b02x02p01n02i02435ent;

ARCHITECTURE c07s03b02x02p01n02i02435arch OF c07s03b02x02p01n02i02435ent IS
  type m1 is array (1 to 3) of integer;
  type m2 is array (1 to 2) of m1;
  constant c: m2 := ((1, 1, 2), (1, 2, 3));  -- No_failure_here
BEGIN
  TESTING: PROCESS
  BEGIN
    assert NOT(c(1)=(1,1,2) and c(2)=(1,2,3))
      report "***PASSED TEST: c07s03b02x02p01n02i02435"
      severity NOTE;
    assert (c(1)=(1,1,2) and c(2)=(1,2,3))
      report "***FAILED TEST: c07s03b02x02p01n02i02435 - Multidimensional aggregates are allowed."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c07s03b02x02p01n02i02435arch;
