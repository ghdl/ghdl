library ieee;use ieee.std_logic_1164;use ieee.numeric_bit_unsigned.all;entity le0el0 is generic(G:integer;G0:integer);port(c:std'l;s:c;--
w:i);end entity le0el0;architecture synthesis of l is
begin
end architecture synthesis;