entity tb is
end tb;

architecture behav of tb is
begin
  p : process
    variable v : natural;
  begin
    v := 5;
    v: null;
  end process;
end behav;
