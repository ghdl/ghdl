use work.a.all;

package b is

  type type_b is record
    something : type_a;
  end record;

end package;
    
