entity repro1 is
  port (a : bit;
        b : bit_vector ());
end repro1;
