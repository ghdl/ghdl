use work.b.all;

package a is

  type type_a is record
    something : type_b;
  end record;

end package;
    
