package n is
function t return n;end;package d is
end;package gen0 is generic(package g is new w generic map(<>));function t return l;end gen0;package body gen0 is use p;function g return l;end gen0;package g is new n;package p is new w generic map(0);architecture beha0 of b is
begin end beha0;