architecture;b';