
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1516.vhd,v 1.2 2001-10-26 16:29:41 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c08s09b00x00p03n01i01516ent IS
END c08s09b00x00p03n01i01516ent;

ARCHITECTURE c08s09b00x00p03n01i01516arch OF c08s09b00x00p03n01i01516ent IS

BEGIN
  TESTING: PROCESS
    type MY_WORD is array (0 to 31) of BIT;
    variable k : integer := 0;
  BEGIN

    for foo in integer range MY_WORD'range loop
      k := k + 1;
    end loop;
    assert NOT(k = 32) 
      report "***PASSED TEST: /c08s09b00x00p03n01i01516"
      severity NOTE;
    assert (k = 32) 
      report "***FAILED TEST: c08s09b00x00p03n01i01516 - FOR loop with a discrete range specification"
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c08s09b00x00p03n01i01516arch;
