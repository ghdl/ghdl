-- comments before design units :p1:
-- :p1: might be multiline
package p1 is
end package;
