entity a is end entity;
architecture b of a is begin end b;
