package function is loop
t((:';