library ieee;
context ieee.ieee_std_context;

entity repro2 is
end repro2; 
