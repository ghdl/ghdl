library ieee;
use ieee.std_logic_1164.all;

library ieee;
use ieee.numeric_std.all;

entity fsm_224 is
	port (
		clock : in  std_logic;
		reset : in  std_logic;
		out40 : out std_logic;
		in2 : in  std_logic;
		in11 : in  std_logic;
		out146 : out std_logic;
		out148 : out std_logic;
		out150 : out std_logic;
		out152 : out std_logic;
		in12 : in  std_logic;
		out153 : out std_logic;
		out154 : out std_logic;
		in13 : in  std_logic;
		out156 : out std_logic;
		out157 : out std_logic;
		out160 : out std_logic;
		out162 : out std_logic;
		out165 : out std_logic;
		out170 : out std_logic;
		out171 : out std_logic;
		out173 : out std_logic;
		out175 : out std_logic;
		out177 : out std_logic;
		out180 : out std_logic;
		out184 : out std_logic;
		in14 : in  std_logic;
		out186 : out std_logic;
		out189 : out std_logic;
		out191 : out std_logic;
		out192 : out std_logic;
		out193 : out std_logic;
		out197 : out std_logic;
		out199 : out std_logic;
		out201 : out std_logic;
		out202 : out std_logic;
		out205 : out std_logic;
		out207 : out std_logic;
		out208 : out std_logic;
		out209 : out std_logic;
		out210 : out std_logic;
		out212 : out std_logic;
		out213 : out std_logic;
		in15 : in  std_logic;
		out221 : out std_logic;
		out222 : out std_logic;
		out224 : out std_logic;
		out225 : out std_logic;
		out228 : out std_logic;
		out229 : out std_logic;
		out230 : out std_logic;
		out231 : out std_logic;
		out99 : out std_logic;
		in6 : in  std_logic;
		out92 : out std_logic;
		out232 : out std_logic;
		in16 : in  std_logic;
		out234 : out std_logic;
		out236 : out std_logic;
		out239 : out std_logic;
		out240 : out std_logic;
		out241 : out std_logic;
		out245 : out std_logic;
		out246 : out std_logic;
		out247 : out std_logic;
		out251 : out std_logic;
		out252 : out std_logic;
		out253 : out std_logic;
		out255 : out std_logic;
		out256 : out std_logic;
		out258 : out std_logic;
		out259 : out std_logic;
		in17 : in  std_logic;
		out263 : out std_logic;
		out264 : out std_logic;
		out266 : out std_logic;
		in18 : in  std_logic;
		out267 : out std_logic;
		out268 : out std_logic;
		out270 : out std_logic;
		out273 : out std_logic;
		out275 : out std_logic;
		out276 : out std_logic;
		in19 : in  std_logic;
		out279 : out std_logic;
		in20 : in  std_logic;
		out281 : out std_logic;
		out282 : out std_logic;
		in21 : in  std_logic;
		out283 : out std_logic;
		out286 : out std_logic;
		out289 : out std_logic;
		out296 : out std_logic;
		out297 : out std_logic;
		out299 : out std_logic;
		out300 : out std_logic;
		out304 : out std_logic;
		out305 : out std_logic;
		in22 : in  std_logic;
		out306 : out std_logic;
		out310 : out std_logic;
		out311 : out std_logic;
		out313 : out std_logic;
		out314 : out std_logic;
		in23 : in  std_logic;
		out316 : out std_logic;
		out317 : out std_logic;
		out320 : out std_logic;
		out322 : out std_logic;
		out324 : out std_logic;
		out325 : out std_logic;
		out326 : out std_logic;
		out328 : out std_logic;
		out332 : out std_logic;
		out333 : out std_logic;
		out334 : out std_logic;
		out335 : out std_logic;
		out338 : out std_logic;
		out339 : out std_logic;
		out341 : out std_logic;
		out342 : out std_logic;
		out344 : out std_logic;
		out93 : out std_logic;
		out98 : out std_logic;
		out85 : out std_logic;
		out87 : out std_logic;
		out88 : out std_logic;
		out80 : out std_logic;
		out82 : out std_logic;
		out83 : out std_logic;
		out84 : out std_logic;
		in5 : in  std_logic;
		out77 : out std_logic;
		out78 : out std_logic;
		out71 : out std_logic;
		out72 : out std_logic;
		in4 : in  std_logic;
		out65 : out std_logic;
		out67 : out std_logic;
		out60 : out std_logic;
		out64 : out std_logic;
		in3 : in  std_logic;
		out59 : out std_logic;
		out53 : out std_logic;
		out55 : out std_logic;
		out49 : out std_logic;
		out44 : out std_logic;
		out104 : out std_logic;
		out107 : out std_logic;
		out111 : out std_logic;
		out112 : out std_logic;
		out114 : out std_logic;
		in7 : in  std_logic;
		out117 : out std_logic;
		out119 : out std_logic;
		out122 : out std_logic;
		in8 : in  std_logic;
		out128 : out std_logic;
		in9 : in  std_logic;
		out129 : out std_logic;
		out130 : out std_logic;
		out133 : out std_logic;
		out134 : out std_logic;
		out136 : out std_logic;
		out137 : out std_logic;
		in10 : in  std_logic;
		out139 : out std_logic;
		out143 : out std_logic;
		out144 : out std_logic;
		out32 : out std_logic;
		out35 : out std_logic;
		out27 : out std_logic;
		out25 : out std_logic;
		out26 : out std_logic;
		in1 : in  std_logic;
		out15 : out std_logic;
		out16 : out std_logic;
		out11 : out std_logic;
		out13 : out std_logic;
		out14 : out std_logic;
		out7 : out std_logic;
		out1 : out std_logic;
		out2 : out std_logic;
		out3 : out std_logic;
		out4 : out std_logic;
		in0 : in  std_logic;
		in24 : in  std_logic;
		out346 : out std_logic;
		out347 : out std_logic;
		out348 : out std_logic;
		out349 : out std_logic;
		in25 : in  std_logic;
		out350 : out std_logic;
		out351 : out std_logic;
		out355 : out std_logic;
		out356 : out std_logic;
		out357 : out std_logic;
		out358 : out std_logic;
		out360 : out std_logic;
		out362 : out std_logic;
		out363 : out std_logic;
		out364 : out std_logic;
		out365 : out std_logic;
		out366 : out std_logic;
		out370 : out std_logic;
		out371 : out std_logic;
		out372 : out std_logic;
		out373 : out std_logic;
		out375 : out std_logic;
		in26 : in  std_logic;
		out376 : out std_logic;
		out378 : out std_logic;
		out379 : out std_logic;
		out381 : out std_logic;
		out382 : out std_logic;
		in27 : in  std_logic;
		out384 : out std_logic;
		in28 : in  std_logic;
		out391 : out std_logic;
		out395 : out std_logic;
		out396 : out std_logic;
		out401 : out std_logic;
		out402 : out std_logic;
		out403 : out std_logic;
		out404 : out std_logic;
		out405 : out std_logic;
		out407 : out std_logic;
		out408 : out std_logic;
		out409 : out std_logic;
		out410 : out std_logic;
		in29 : in  std_logic;
		out412 : out std_logic;
		out414 : out std_logic;
		out415 : out std_logic;
		out417 : out std_logic;
		out418 : out std_logic;
		out419 : out std_logic;
		out420 : out std_logic;
		out422 : out std_logic;
		out424 : out std_logic;
		out425 : out std_logic;
		out426 : out std_logic;
		in30 : in  std_logic;
		out428 : out std_logic;
		out429 : out std_logic;
		out432 : out std_logic;
		out433 : out std_logic;
		out434 : out std_logic;
		out437 : out std_logic;
		out440 : out std_logic;
		out441 : out std_logic;
		in31 : in  std_logic;
		out443 : out std_logic;
		in32 : in  std_logic;
		out445 : out std_logic;
		out447 : out std_logic;
		out448 : out std_logic;
		out450 : out std_logic;
		in33 : in  std_logic;
		out453 : out std_logic;
		out455 : out std_logic;
		out458 : out std_logic;
		in34 : in  std_logic;
		out462 : out std_logic;
		out464 : out std_logic;
		out467 : out std_logic;
		out468 : out std_logic;
		out472 : out std_logic;
		in35 : in  std_logic;
		out478 : out std_logic;
		out479 : out std_logic;
		out480 : out std_logic;
		out487 : out std_logic;
		out488 : out std_logic;
		in36 : in  std_logic;
		out491 : out std_logic;
		out496 : out std_logic;
		out497 : out std_logic;
		out498 : out std_logic;
		out500 : out std_logic;
		out504 : out std_logic;
		out505 : out std_logic;
		in37 : in  std_logic;
		out506 : out std_logic;
		out508 : out std_logic;
		in38 : in  std_logic;
		out510 : out std_logic;
		out513 : out std_logic;
		out514 : out std_logic;
		out515 : out std_logic;
		out517 : out std_logic;
		out519 : out std_logic;
		in39 : in  std_logic;
		out523 : out std_logic;
		out526 : out std_logic;
		out527 : out std_logic;
		out528 : out std_logic;
		out530 : out std_logic;
		out531 : out std_logic;
		out533 : out std_logic;
		out534 : out std_logic;
		out537 : out std_logic;
		out538 : out std_logic;
		out549 : out std_logic;
		out558 : out std_logic;
		out559 : out std_logic;
		out561 : out std_logic;
		in40 : in  std_logic;
		out566 : out std_logic;
		out567 : out std_logic;
		out568 : out std_logic;
		out569 : out std_logic;
		out570 : out std_logic;
		out572 : out std_logic;
		out574 : out std_logic;
		out575 : out std_logic;
		out577 : out std_logic;
		in41 : in  std_logic;
		out578 : out std_logic;
		out581 : out std_logic;
		out589 : out std_logic;
		out590 : out std_logic;
		out595 : out std_logic;
		out597 : out std_logic;
		out599 : out std_logic;
		out601 : out std_logic;
		out602 : out std_logic;
		out607 : out std_logic;
		out610 : out std_logic;
		out612 : out std_logic;
		in42 : in  std_logic;
		out614 : out std_logic;
		out621 : out std_logic;
		out628 : out std_logic;
		out635 : out std_logic;
		out636 : out std_logic;
		out638 : out std_logic;
		out640 : out std_logic;
		out643 : out std_logic;
		out646 : out std_logic;
		out649 : out std_logic;
		out651 : out std_logic;
		out656 : out std_logic;
		in43 : in  std_logic;
		out658 : out std_logic;
		out659 : out std_logic;
		out661 : out std_logic;
		out663 : out std_logic;
		out664 : out std_logic;
		in44 : in  std_logic;
		out667 : out std_logic;
		out668 : out std_logic;
		out670 : out std_logic;
		out672 : out std_logic;
		out674 : out std_logic;
		in45 : in  std_logic;
		out679 : out std_logic;
		out681 : out std_logic;
		out683 : out std_logic;
		out686 : out std_logic;
		out688 : out std_logic;
		out690 : out std_logic;
		out692 : out std_logic;
		out694 : out std_logic;
		out696 : out std_logic;
		out697 : out std_logic;
		out698 : out std_logic;
		out699 : out std_logic;
		out700 : out std_logic;
		out703 : out std_logic;
		out704 : out std_logic;
		out706 : out std_logic;
		out708 : out std_logic;
		out710 : out std_logic;
		out712 : out std_logic;
		out715 : out std_logic;
		out718 : out std_logic;
		in46 : in  std_logic;
		out722 : out std_logic;
		out724 : out std_logic;
		out726 : out std_logic;
		out728 : out std_logic;
		out731 : out std_logic;
		out733 : out std_logic;
		out734 : out std_logic;
		out737 : out std_logic;
		out739 : out std_logic;
		out740 : out std_logic;
		out743 : out std_logic;
		out745 : out std_logic;
		out746 : out std_logic;
		in47 : in  std_logic;
		out749 : out std_logic;
		out753 : out std_logic;
		out755 : out std_logic;
		out759 : out std_logic;
		in48 : in  std_logic;
		out762 : out std_logic;
		out764 : out std_logic;
		out765 : out std_logic;
		out767 : out std_logic;
		out768 : out std_logic;
		in49 : in  std_logic;
		out772 : out std_logic;
		in50 : in  std_logic;
		out775 : out std_logic;
		out776 : out std_logic;
		out778 : out std_logic;
		out783 : out std_logic;
		out784 : out std_logic;
		out787 : out std_logic;
		out791 : out std_logic;
		in51 : in  std_logic;
		out794 : out std_logic;
		out795 : out std_logic;
		in52 : in  std_logic;
		out799 : out std_logic;
		out802 : out std_logic;
		out806 : out std_logic;
		out809 : out std_logic;
		out812 : out std_logic;
		out815 : out std_logic;
		out826 : out std_logic;
		out828 : out std_logic;
		in53 : in  std_logic;
		in54 : in  std_logic;
		out843 : out std_logic;
		out848 : out std_logic;
		out852 : out std_logic;
		in55 : in  std_logic;
		out855 : out std_logic;
		out858 : out std_logic;
		in56 : in  std_logic;
		out860 : out std_logic;
		out861 : out std_logic;
		out863 : out std_logic;
		out866 : out std_logic;
		out872 : out std_logic;
		in57 : in  std_logic;
		out874 : out std_logic;
		out876 : out std_logic;
		out879 : out std_logic;
		out882 : out std_logic;
		out886 : out std_logic;
		out887 : out std_logic;
		in58 : in  std_logic;
		out888 : out std_logic;
		out892 : out std_logic;
		out894 : out std_logic;
		out895 : out std_logic;
		out896 : out std_logic;
		out901 : out std_logic;
		out902 : out std_logic;
		out903 : out std_logic;
		out905 : out std_logic;
		out907 : out std_logic;
		out918 : out std_logic;
		out920 : out std_logic;
		out921 : out std_logic;
		out923 : out std_logic;
		out925 : out std_logic;
		out928 : out std_logic;
		out929 : out std_logic;
		out931 : out std_logic;
		out933 : out std_logic;
		out936 : out std_logic;
		out937 : out std_logic;
		out938 : out std_logic;
		out939 : out std_logic;
		out942 : out std_logic;
		out943 : out std_logic;
		out944 : out std_logic;
		out947 : out std_logic;
		out948 : out std_logic;
		out949 : out std_logic;
		out951 : out std_logic;
		in59 : in  std_logic;
		out952 : out std_logic;
		out953 : out std_logic;
		out955 : out std_logic;
		out956 : out std_logic;
		out957 : out std_logic;
		out958 : out std_logic;
		in60 : in  std_logic;
		in61 : in  std_logic;
		out962 : out std_logic;
		out963 : out std_logic;
		out972 : out std_logic;
		out973 : out std_logic;
		out974 : out std_logic;
		in62 : in  std_logic;
		out978 : out std_logic;
		out979 : out std_logic;
		out981 : out std_logic;
		out982 : out std_logic;
		out985 : out std_logic;
		out986 : out std_logic;
		out989 : out std_logic;
		in63 : in  std_logic;
		in64 : in  std_logic;
		in65 : in  std_logic;
		in66 : in  std_logic;
		in67 : in  std_logic;
		in68 : in  std_logic;
		in69 : in  std_logic;
		in70 : in  std_logic;
		in71 : in  std_logic;
		in72 : in  std_logic;
		in73 : in  std_logic;
		in74 : in  std_logic;
		in75 : in  std_logic;
		in76 : in  std_logic;
		in77 : in  std_logic;
		in78 : in  std_logic;
		out990 : out std_logic;
		out991 : out std_logic;
		out993 : out std_logic;
		out994 : out std_logic;
		out996 : out std_logic;
		out997 : out std_logic;
		out998 : out std_logic;
		out999 : out std_logic;
		out1000 : out std_logic;
		out1002 : out std_logic;
		out1003 : out std_logic;
		out1005 : out std_logic;
		out1006 : out std_logic;
		out1007 : out std_logic;
		out1009 : out std_logic;
		out1011 : out std_logic;
		out1012 : out std_logic;
		out1013 : out std_logic;
		out1014 : out std_logic;
		out1015 : out std_logic;
		out1016 : out std_logic;
		out1018 : out std_logic;
		out1019 : out std_logic;
		out1021 : out std_logic;
		out1022 : out std_logic;
		out1024 : out std_logic;
		out1026 : out std_logic;
		out1027 : out std_logic;
		out1029 : out std_logic;
		out1030 : out std_logic;
		out1032 : out std_logic;
		out1033 : out std_logic;
		out1035 : out std_logic;
		out1036 : out std_logic;
		out1037 : out std_logic;
		out1057 : out std_logic;
		out1068 : out std_logic;
		out1069 : out std_logic;
		out1070 : out std_logic;
		out1072 : out std_logic;
		out1073 : out std_logic;
		out1075 : out std_logic;
		out1078 : out std_logic;
		out1080 : out std_logic;
		out1082 : out std_logic;
		out1083 : out std_logic;
		out1084 : out std_logic;
		out1085 : out std_logic;
		out1088 : out std_logic;
		out1089 : out std_logic;
		out1091 : out std_logic;
		out1092 : out std_logic;
		out1094 : out std_logic;
		out1096 : out std_logic;
		out1098 : out std_logic;
		out1101 : out std_logic;
		out1104 : out std_logic;
		out1107 : out std_logic;
		out1109 : out std_logic;
		out1111 : out std_logic;
		out1114 : out std_logic;
		out1119 : out std_logic;
		out1121 : out std_logic;
		out1125 : out std_logic;
		out1126 : out std_logic;
		out1128 : out std_logic;
		out1131 : out std_logic;
		out1134 : out std_logic;
		out1137 : out std_logic;
		out1139 : out std_logic;
		out1141 : out std_logic;
		out1145 : out std_logic;
		out1146 : out std_logic;
		out1147 : out std_logic;
		out1150 : out std_logic;
		out1151 : out std_logic;
		out1152 : out std_logic;
		out1155 : out std_logic;
		out1158 : out std_logic;
		out1160 : out std_logic;
		out1164 : out std_logic;
		out1166 : out std_logic;
		out1169 : out std_logic;
		out1171 : out std_logic;
		out1174 : out std_logic;
		out1175 : out std_logic;
		out1176 : out std_logic;
		out1180 : out std_logic;
		out1181 : out std_logic;
		out1182 : out std_logic;
		out1185 : out std_logic;
		out1186 : out std_logic;
		out1187 : out std_logic;
		out1190 : out std_logic;
		out1213 : out std_logic;
		out1215 : out std_logic;
		out1217 : out std_logic;
		out1220 : out std_logic;
		out1221 : out std_logic;
		out1223 : out std_logic;
		out1228 : out std_logic;
		out1229 : out std_logic;
		out1231 : out std_logic;
		out1235 : out std_logic;
		out1236 : out std_logic;
		out1240 : out std_logic;
		out1243 : out std_logic;
		out1250 : out std_logic;
		out1252 : out std_logic;
		out1253 : out std_logic;
		out1258 : out std_logic;
		out1262 : out std_logic;
		out1266 : out std_logic;
		out1269 : out std_logic;
		out1275 : out std_logic;
		out1278 : out std_logic;
		out1279 : out std_logic;
		out1284 : out std_logic;
		out1286 : out std_logic;
		out1287 : out std_logic;
		out1289 : out std_logic;
		out1290 : out std_logic;
		out1292 : out std_logic;
		out1293 : out std_logic;
		out1295 : out std_logic;
		out1298 : out std_logic;
		out1301 : out std_logic;
		out1302 : out std_logic;
		out1303 : out std_logic;
		out1308 : out std_logic;
		out1309 : out std_logic;
		out1311 : out std_logic;
		out1318 : out std_logic;
		out1319 : out std_logic;
		out1320 : out std_logic;
		out1323 : out std_logic;
		out1324 : out std_logic;
		out1326 : out std_logic;
		out1327 : out std_logic;
		out1329 : out std_logic;
		out1337 : out std_logic;
		out1339 : out std_logic;
		out1340 : out std_logic;
		out1341 : out std_logic;
		out1344 : out std_logic;
		out1346 : out std_logic;
		out1349 : out std_logic;
		out1353 : out std_logic;
		out1356 : out std_logic;
		out1362 : out std_logic;
		out1363 : out std_logic;
		out1364 : out std_logic;
		out1365 : out std_logic;
		out1366 : out std_logic;
		out1368 : out std_logic;
		out1370 : out std_logic;
		out1375 : out std_logic;
		out1378 : out std_logic;
		out1381 : out std_logic;
		out1383 : out std_logic;
		out1387 : out std_logic
	);
end fsm_224;

architecture augh of fsm_224 is

	signal state_cur  : std_logic_vector(0 to 473) := (457 => '1', others => '0');
	signal state_next : std_logic_vector(0 to 473) := (457 => '1', others => '0');

	-- Buffers for outputs
	signal out1057_buf : std_logic := '0';
	signal out1057_bufn : std_logic;
	signal out59_buf : std_logic := '0';
	signal out59_bufn : std_logic;
	signal out447_buf : std_logic := '0';
	signal out447_bufn : std_logic;
	signal out157_buf : std_logic := '0';
	signal out157_bufn : std_logic;
	signal out450_buf : std_logic := '0';
	signal out450_bufn : std_logic;
	signal out1012_buf : std_logic := '0';
	signal out1012_bufn : std_logic;
	signal out1072_buf : std_logic := '0';
	signal out1072_bufn : std_logic;
	signal out999_buf : std_logic := '0';
	signal out999_bufn : std_logic;
	signal out437_buf : std_logic := '0';
	signal out437_bufn : std_logic;
	signal out415_buf : std_logic := '0';
	signal out415_bufn : std_logic;
	signal out426_buf : std_logic := '0';
	signal out426_bufn : std_logic;
	signal out375_buf : std_logic := '0';
	signal out375_bufn : std_logic;
	signal out704_buf : std_logic := '0';
	signal out704_bufn : std_logic;
	signal out973_buf : std_logic := '0';
	signal out973_bufn : std_logic;
	signal out11_buf : std_logic := '0';
	signal out11_bufn : std_logic;
	signal out549_buf : std_logic := '0';
	signal out549_bufn : std_logic;
	signal out453_buf : std_logic := '0';
	signal out453_bufn : std_logic;
	signal out1231_buf : std_logic := '0';
	signal out1231_bufn : std_logic;
	signal out87_buf : std_logic := '0';
	signal out87_bufn : std_logic;
	signal out401_buf : std_logic := '0';
	signal out401_bufn : std_logic;
	signal out990_buf : std_logic := '0';
	signal out990_bufn : std_logic;
	signal out378_buf : std_logic := '0';
	signal out378_bufn : std_logic;
	signal out1302_buf : std_logic := '0';
	signal out1302_bufn : std_logic;
	signal out27_buf : std_logic := '0';
	signal out27_bufn : std_logic;
	signal out569_buf : std_logic := '0';
	signal out569_bufn : std_logic;
	signal out1030_buf : std_logic := '0';
	signal out1030_bufn : std_logic;
	signal out537_buf : std_logic := '0';
	signal out537_bufn : std_logic;
	signal out77_buf : std_logic := '0';
	signal out77_bufn : std_logic;
	signal out1318_buf : std_logic := '0';
	signal out1318_bufn : std_logic;
	signal out533_buf : std_logic := '0';
	signal out533_bufn : std_logic;
	signal out32_buf : std_logic := '0';
	signal out32_bufn : std_logic;
	signal out1027_buf : std_logic := '0';
	signal out1027_bufn : std_logic;
	signal out599_buf : std_logic := '0';
	signal out599_bufn : std_logic;
	signal out668_buf : std_logic := '0';
	signal out668_bufn : std_logic;
	signal out568_buf : std_logic := '0';
	signal out568_bufn : std_logic;
	signal out225_buf : std_logic := '0';
	signal out225_bufn : std_logic;
	signal out700_buf : std_logic := '0';
	signal out700_bufn : std_logic;
	signal out638_buf : std_logic := '0';
	signal out638_bufn : std_logic;
	signal out670_buf : std_logic := '0';
	signal out670_bufn : std_logic;
	signal out433_buf : std_logic := '0';
	signal out433_bufn : std_logic;
	signal out896_buf : std_logic := '0';
	signal out896_bufn : std_logic;
	signal out575_buf : std_logic := '0';
	signal out575_bufn : std_logic;
	signal out428_buf : std_logic := '0';
	signal out428_bufn : std_logic;
	signal out72_buf : std_logic := '0';
	signal out72_bufn : std_logic;
	signal out404_buf : std_logic := '0';
	signal out404_bufn : std_logic;
	signal out98_buf : std_logic := '0';
	signal out98_bufn : std_logic;
	signal out67_buf : std_logic := '0';
	signal out67_bufn : std_logic;
	signal out635_buf : std_logic := '0';
	signal out635_bufn : std_logic;
	signal out381_buf : std_logic := '0';
	signal out381_bufn : std_logic;
	signal out222_buf : std_logic := '0';
	signal out222_bufn : std_logic;
	signal out339_buf : std_logic := '0';
	signal out339_bufn : std_logic;
	signal out268_buf : std_logic := '0';
	signal out268_bufn : std_logic;
	signal out419_buf : std_logic := '0';
	signal out419_bufn : std_logic;
	signal out559_buf : std_logic := '0';
	signal out559_bufn : std_logic;
	signal out1002_buf : std_logic := '0';
	signal out1002_bufn : std_logic;
	signal out1006_buf : std_logic := '0';
	signal out1006_bufn : std_logic;
	signal out276_buf : std_logic := '0';
	signal out276_bufn : std_logic;
	signal out205_buf : std_logic := '0';
	signal out205_bufn : std_logic;
	signal out943_buf : std_logic := '0';
	signal out943_bufn : std_logic;
	signal out1080_buf : std_logic := '0';
	signal out1080_bufn : std_logic;
	signal out408_buf : std_logic := '0';
	signal out408_bufn : std_logic;
	signal out252_buf : std_logic := '0';
	signal out252_bufn : std_logic;
	signal out71_buf : std_logic := '0';
	signal out71_bufn : std_logic;
	signal out672_buf : std_logic := '0';
	signal out672_bufn : std_logic;
	signal out357_buf : std_logic := '0';
	signal out357_bufn : std_logic;
	signal out441_buf : std_logic := '0';
	signal out441_bufn : std_logic;
	signal out1084_buf : std_logic := '0';
	signal out1084_bufn : std_logic;
	signal out144_buf : std_logic := '0';
	signal out144_bufn : std_logic;
	signal out574_buf : std_logic := '0';
	signal out574_bufn : std_logic;
	signal out210_buf : std_logic := '0';
	signal out210_bufn : std_logic;
	signal out128_buf : std_logic := '0';
	signal out128_bufn : std_logic;
	signal out360_buf : std_logic := '0';
	signal out360_bufn : std_logic;
	signal out948_buf : std_logic := '0';
	signal out948_bufn : std_logic;
	signal out506_buf : std_logic := '0';
	signal out506_bufn : std_logic;
	signal out207_buf : std_logic := '0';
	signal out207_bufn : std_logic;
	signal out1083_buf : std_logic := '0';
	signal out1083_bufn : std_logic;
	signal out491_buf : std_logic := '0';
	signal out491_bufn : std_logic;
	signal out4_buf : std_logic := '0';
	signal out4_bufn : std_logic;
	signal out784_buf : std_logic := '0';
	signal out784_bufn : std_logic;
	signal out3_buf : std_logic := '0';
	signal out3_bufn : std_logic;
	signal out746_buf : std_logic := '0';
	signal out746_bufn : std_logic;
	signal out528_buf : std_logic := '0';
	signal out528_bufn : std_logic;
	signal out372_buf : std_logic := '0';
	signal out372_bufn : std_logic;
	signal out418_buf : std_logic := '0';
	signal out418_bufn : std_logic;
	signal out708_buf : std_logic := '0';
	signal out708_bufn : std_logic;
	signal out706_buf : std_logic := '0';
	signal out706_bufn : std_logic;
	signal out445_buf : std_logic := '0';
	signal out445_bufn : std_logic;
	signal out1021_buf : std_logic := '0';
	signal out1021_bufn : std_logic;
	signal out405_buf : std_logic := '0';
	signal out405_bufn : std_logic;
	signal out764_buf : std_logic := '0';
	signal out764_bufn : std_logic;
	signal out581_buf : std_logic := '0';
	signal out581_bufn : std_logic;
	signal out776_buf : std_logic := '0';
	signal out776_bufn : std_logic;
	signal out213_buf : std_logic := '0';
	signal out213_bufn : std_logic;
	signal out674_buf : std_logic := '0';
	signal out674_bufn : std_logic;
	signal out1326_buf : std_logic := '0';
	signal out1326_bufn : std_logic;
	signal out334_buf : std_logic := '0';
	signal out334_bufn : std_logic;
	signal out843_buf : std_logic := '0';
	signal out843_bufn : std_logic;
	signal out175_buf : std_logic := '0';
	signal out175_bufn : std_logic;
	signal out1036_buf : std_logic := '0';
	signal out1036_bufn : std_logic;
	signal out1015_buf : std_logic := '0';
	signal out1015_bufn : std_logic;
	signal out236_buf : std_logic := '0';
	signal out236_bufn : std_logic;
	signal out395_buf : std_logic := '0';
	signal out395_bufn : std_logic;
	signal out1340_buf : std_logic := '0';
	signal out1340_bufn : std_logic;
	signal out993_buf : std_logic := '0';
	signal out993_bufn : std_logic;
	signal out356_buf : std_logic := '0';
	signal out356_bufn : std_logic;
	signal out273_buf : std_logic := '0';
	signal out273_bufn : std_logic;
	signal out403_buf : std_logic := '0';
	signal out403_bufn : std_logic;
	signal out286_buf : std_logic := '0';
	signal out286_bufn : std_logic;
	signal out364_buf : std_logic := '0';
	signal out364_bufn : std_logic;
	signal out697_buf : std_logic := '0';
	signal out697_bufn : std_logic;
	signal out283_buf : std_logic := '0';
	signal out283_bufn : std_logic;
	signal out282_buf : std_logic := '0';
	signal out282_bufn : std_logic;
	signal out1319_buf : std_logic := '0';
	signal out1319_bufn : std_logic;
	signal out409_buf : std_logic := '0';
	signal out409_bufn : std_logic;
	signal out1092_buf : std_logic := '0';
	signal out1092_bufn : std_logic;
	signal out1075_buf : std_logic := '0';
	signal out1075_bufn : std_logic;
	signal out925_buf : std_logic := '0';
	signal out925_bufn : std_logic;
	signal out78_buf : std_logic := '0';
	signal out78_bufn : std_logic;
	signal out1089_buf : std_logic := '0';
	signal out1089_bufn : std_logic;
	signal out362_buf : std_logic := '0';
	signal out362_bufn : std_logic;
	signal out982_buf : std_logic := '0';
	signal out982_bufn : std_logic;
	signal out979_buf : std_logic := '0';
	signal out979_bufn : std_logic;
	signal out952_buf : std_logic := '0';
	signal out952_bufn : std_logic;
	signal out1109_buf : std_logic := '0';
	signal out1109_bufn : std_logic;
	signal out16_buf : std_logic := '0';
	signal out16_bufn : std_logic;
	signal out703_buf : std_logic := '0';
	signal out703_bufn : std_logic;
	signal out371_buf : std_logic := '0';
	signal out371_bufn : std_logic;
	signal out956_buf : std_logic := '0';
	signal out956_bufn : std_logic;
	signal out1107_buf : std_logic := '0';
	signal out1107_bufn : std_logic;
	signal out1033_buf : std_logic := '0';
	signal out1033_bufn : std_logic;
	signal out148_buf : std_logic := '0';
	signal out148_bufn : std_logic;
	signal out351_buf : std_logic := '0';
	signal out351_bufn : std_logic;
	signal out740_buf : std_logic := '0';
	signal out740_bufn : std_logic;
	signal out391_buf : std_logic := '0';
	signal out391_bufn : std_logic;
	signal out129_buf : std_logic := '0';
	signal out129_bufn : std_logic;
	signal out338_buf : std_logic := '0';
	signal out338_bufn : std_logic;
	signal out425_buf : std_logic := '0';
	signal out425_bufn : std_logic;
	signal out1078_buf : std_logic := '0';
	signal out1078_bufn : std_logic;
	signal out349_buf : std_logic := '0';
	signal out349_bufn : std_logic;
	signal out590_buf : std_logic := '0';
	signal out590_bufn : std_logic;
	signal out325_buf : std_logic := '0';
	signal out325_bufn : std_logic;
	signal out112_buf : std_logic := '0';
	signal out112_bufn : std_logic;
	signal out224_buf : std_logic := '0';
	signal out224_bufn : std_logic;
	signal out1220_buf : std_logic := '0';
	signal out1220_bufn : std_logic;
	signal out1250_buf : std_logic := '0';
	signal out1250_bufn : std_logic;
	signal out365_buf : std_logic := '0';
	signal out365_bufn : std_logic;
	signal out699_buf : std_logic := '0';
	signal out699_bufn : std_logic;
	signal out488_buf : std_logic := '0';
	signal out488_bufn : std_logic;
	signal out1069_buf : std_logic := '0';
	signal out1069_bufn : std_logic;
	signal out530_buf : std_logic := '0';
	signal out530_bufn : std_logic;
	signal out326_buf : std_logic := '0';
	signal out326_bufn : std_logic;
	signal out602_buf : std_logic := '0';
	signal out602_bufn : std_logic;
	signal out83_buf : std_logic := '0';
	signal out83_bufn : std_logic;
	signal out311_buf : std_logic := '0';
	signal out311_bufn : std_logic;
	signal out253_buf : std_logic := '0';
	signal out253_bufn : std_logic;
	signal out209_buf : std_logic := '0';
	signal out209_bufn : std_logic;
	signal out1240_buf : std_logic := '0';
	signal out1240_bufn : std_logic;
	signal out1018_buf : std_logic := '0';
	signal out1018_bufn : std_logic;
	signal out1152_buf : std_logic := '0';
	signal out1152_bufn : std_logic;
	signal out1236_buf : std_logic := '0';
	signal out1236_bufn : std_logic;
	signal out130_buf : std_logic := '0';
	signal out130_bufn : std_logic;
	signal out567_buf : std_logic := '0';
	signal out567_bufn : std_logic;
	signal out646_buf : std_logic := '0';
	signal out646_bufn : std_logic;

	-- Function calls: return IDs
	signal funccall0 : natural range 0 to 18 := 0;
	signal funccall0_next : natural range 0 to 18 := 0;
	signal funccall1 : natural range 0 to 6 := 0;
	signal funccall1_next : natural range 0 to 6 := 0;
	signal funccall2 : natural range 0 to 2 := 0;
	signal funccall2_next : natural range 0 to 2 := 0;
	signal funccall3 : natural range 0 to 3 := 0;
	signal funccall3_next : natural range 0 to 3 := 0;
	signal funccall4 : natural range 0 to 1 := 0;
	signal funccall4_next : natural range 0 to 1 := 0;
	signal funccall5 : natural range 0 to 1 := 0;
	signal funccall5_next : natural range 0 to 1 := 0;
	signal funccall6 : natural range 0 to 1 := 0;
	signal funccall6_next : natural range 0 to 1 := 0;
	signal funccall7 : natural range 0 to 4 := 0;
	signal funccall7_next : natural range 0 to 4 := 0;
	signal funccall8 : natural range 0 to 1 := 0;
	signal funccall8_next : natural range 0 to 1 := 0;
	signal funccall9 : natural range 0 to 3 := 0;
	signal funccall9_next : natural range 0 to 3 := 0;

	-- A utility function to convert bool to std_logic
	function to_stdl (b: boolean) return std_logic is
	begin
		if b = true then
			return '1';
		end if;
		return '0';
	end function;

begin

	-- Sequential process
	-- Set the current state

	process (clock)
	begin
		if rising_edge(clock) then

			-- Next state
			state_cur <= state_next;
			-- Buffers for outputs
			out1057_buf <= out1057_bufn;
			out59_buf <= out59_bufn;
			out447_buf <= out447_bufn;
			out157_buf <= out157_bufn;
			out450_buf <= out450_bufn;
			out1012_buf <= out1012_bufn;
			out1072_buf <= out1072_bufn;
			out999_buf <= out999_bufn;
			out437_buf <= out437_bufn;
			out415_buf <= out415_bufn;
			out426_buf <= out426_bufn;
			out375_buf <= out375_bufn;
			out704_buf <= out704_bufn;
			out973_buf <= out973_bufn;
			out11_buf <= out11_bufn;
			out549_buf <= out549_bufn;
			out453_buf <= out453_bufn;
			out1231_buf <= out1231_bufn;
			out87_buf <= out87_bufn;
			out401_buf <= out401_bufn;
			out990_buf <= out990_bufn;
			out378_buf <= out378_bufn;
			out1302_buf <= out1302_bufn;
			out27_buf <= out27_bufn;
			out569_buf <= out569_bufn;
			out1030_buf <= out1030_bufn;
			out537_buf <= out537_bufn;
			out77_buf <= out77_bufn;
			out1318_buf <= out1318_bufn;
			out533_buf <= out533_bufn;
			out32_buf <= out32_bufn;
			out1027_buf <= out1027_bufn;
			out599_buf <= out599_bufn;
			out668_buf <= out668_bufn;
			out568_buf <= out568_bufn;
			out225_buf <= out225_bufn;
			out700_buf <= out700_bufn;
			out638_buf <= out638_bufn;
			out670_buf <= out670_bufn;
			out433_buf <= out433_bufn;
			out896_buf <= out896_bufn;
			out575_buf <= out575_bufn;
			out428_buf <= out428_bufn;
			out72_buf <= out72_bufn;
			out404_buf <= out404_bufn;
			out98_buf <= out98_bufn;
			out67_buf <= out67_bufn;
			out635_buf <= out635_bufn;
			out381_buf <= out381_bufn;
			out222_buf <= out222_bufn;
			out339_buf <= out339_bufn;
			out268_buf <= out268_bufn;
			out419_buf <= out419_bufn;
			out559_buf <= out559_bufn;
			out1002_buf <= out1002_bufn;
			out1006_buf <= out1006_bufn;
			out276_buf <= out276_bufn;
			out205_buf <= out205_bufn;
			out943_buf <= out943_bufn;
			out1080_buf <= out1080_bufn;
			out408_buf <= out408_bufn;
			out252_buf <= out252_bufn;
			out71_buf <= out71_bufn;
			out672_buf <= out672_bufn;
			out357_buf <= out357_bufn;
			out441_buf <= out441_bufn;
			out1084_buf <= out1084_bufn;
			out144_buf <= out144_bufn;
			out574_buf <= out574_bufn;
			out210_buf <= out210_bufn;
			out128_buf <= out128_bufn;
			out360_buf <= out360_bufn;
			out948_buf <= out948_bufn;
			out506_buf <= out506_bufn;
			out207_buf <= out207_bufn;
			out1083_buf <= out1083_bufn;
			out491_buf <= out491_bufn;
			out4_buf <= out4_bufn;
			out784_buf <= out784_bufn;
			out3_buf <= out3_bufn;
			out746_buf <= out746_bufn;
			out528_buf <= out528_bufn;
			out372_buf <= out372_bufn;
			out418_buf <= out418_bufn;
			out708_buf <= out708_bufn;
			out706_buf <= out706_bufn;
			out445_buf <= out445_bufn;
			out1021_buf <= out1021_bufn;
			out405_buf <= out405_bufn;
			out764_buf <= out764_bufn;
			out581_buf <= out581_bufn;
			out776_buf <= out776_bufn;
			out213_buf <= out213_bufn;
			out674_buf <= out674_bufn;
			out1326_buf <= out1326_bufn;
			out334_buf <= out334_bufn;
			out843_buf <= out843_bufn;
			out175_buf <= out175_bufn;
			out1036_buf <= out1036_bufn;
			out1015_buf <= out1015_bufn;
			out236_buf <= out236_bufn;
			out395_buf <= out395_bufn;
			out1340_buf <= out1340_bufn;
			out993_buf <= out993_bufn;
			out356_buf <= out356_bufn;
			out273_buf <= out273_bufn;
			out403_buf <= out403_bufn;
			out286_buf <= out286_bufn;
			out364_buf <= out364_bufn;
			out697_buf <= out697_bufn;
			out283_buf <= out283_bufn;
			out282_buf <= out282_bufn;
			out1319_buf <= out1319_bufn;
			out409_buf <= out409_bufn;
			out1092_buf <= out1092_bufn;
			out1075_buf <= out1075_bufn;
			out925_buf <= out925_bufn;
			out78_buf <= out78_bufn;
			out1089_buf <= out1089_bufn;
			out362_buf <= out362_bufn;
			out982_buf <= out982_bufn;
			out979_buf <= out979_bufn;
			out952_buf <= out952_bufn;
			out1109_buf <= out1109_bufn;
			out16_buf <= out16_bufn;
			out703_buf <= out703_bufn;
			out371_buf <= out371_bufn;
			out956_buf <= out956_bufn;
			out1107_buf <= out1107_bufn;
			out1033_buf <= out1033_bufn;
			out148_buf <= out148_bufn;
			out351_buf <= out351_bufn;
			out740_buf <= out740_bufn;
			out391_buf <= out391_bufn;
			out129_buf <= out129_bufn;
			out338_buf <= out338_bufn;
			out425_buf <= out425_bufn;
			out1078_buf <= out1078_bufn;
			out349_buf <= out349_bufn;
			out590_buf <= out590_bufn;
			out325_buf <= out325_bufn;
			out112_buf <= out112_bufn;
			out224_buf <= out224_bufn;
			out1220_buf <= out1220_bufn;
			out1250_buf <= out1250_bufn;
			out365_buf <= out365_bufn;
			out699_buf <= out699_bufn;
			out488_buf <= out488_bufn;
			out1069_buf <= out1069_bufn;
			out530_buf <= out530_bufn;
			out326_buf <= out326_bufn;
			out602_buf <= out602_bufn;
			out83_buf <= out83_bufn;
			out311_buf <= out311_bufn;
			out253_buf <= out253_bufn;
			out209_buf <= out209_bufn;
			out1240_buf <= out1240_bufn;
			out1018_buf <= out1018_bufn;
			out1152_buf <= out1152_bufn;
			out1236_buf <= out1236_bufn;
			out130_buf <= out130_bufn;
			out567_buf <= out567_bufn;
			out646_buf <= out646_bufn;
			-- Function calls: return IDs
			funccall0 <= funccall0_next;
			funccall1 <= funccall1_next;
			funccall2 <= funccall2_next;
			funccall3 <= funccall3_next;
			funccall4 <= funccall4_next;
			funccall5 <= funccall5_next;
			funccall6 <= funccall6_next;
			funccall7 <= funccall7_next;
			funccall8 <= funccall8_next;
			funccall9 <= funccall9_next;

		end if;
	end process;

	-- Function calls: The call IDs

	-- Function 'read_byte'
	funccall0_next <=
		0 when ( state_cur(130) and in33 ) = '1' else
		2 when ( state_cur(130) and not ( in33 ) ) = '1' else
		18 when ( state_cur(137) and not ( in34 ) ) = '1' else
		17 when ( state_cur(148) and in36 ) = '1' else
		16 when ( state_cur(160) and in38 ) = '1' else
		15 when ( state_cur(170) and in39 ) = '1' else
		14 when ( state_cur(179) and in40 ) = '1' else
		10 when ( state_cur(207) and to_stdl(funccall1 = 3) ) = '1' else
		5 when ( state_cur(207) and to_stdl(funccall1 = 0) ) = '1' else
		12 when state_cur(211) = '1' else
		11 when ( state_cur(212) and in43 ) = '1' else
		9 when state_cur(237) = '1' else
		8 when state_cur(238) = '1' else
		7 when state_cur(242) = '1' else
		6 when state_cur(243) = '1' else
		2 when ( state_cur(246) and not ( in46 ) ) = '1' else
		3 when ( state_cur(249) and in47 ) = '1' else
		4 when ( state_cur(249) and not ( in47 ) ) = '1' else
		4 when ( state_cur(251) and in48 ) = '1' else
		13 when ( state_cur(338) and in52 ) = '1' else
		1 when ( state_cur(396) and to_stdl(funccall0 = 0) ) = '1' else
		funccall0;
	-- Function 'read_word'
	funccall1_next <=
		5 when ( state_cur(126) and not ( in32 ) and in31 ) = '1' else
		4 when ( state_cur(126) and not ( in32 ) and not ( in31 ) and in30 ) = '1' else
		3 when ( state_cur(126) and not ( in32 ) and not ( in31 ) and not ( in30 ) and in29 ) = '1' else
		0 when ( state_cur(126) and not ( in32 ) and not ( in31 ) and not ( in30 ) and not ( in29 ) and in28 ) = '1' else
		6 when ( state_cur(137) and in34 ) = '1' else
		2 when state_cur(244) = '1' else
		1 when ( state_cur(396) and to_stdl(funccall0 = 5) ) = '1' else
		funccall1;
	-- Function 'pgetc'
	funccall2_next <=
		1 when state_cur(72) = '1' else
		2 when ( state_cur(73) and not ( in20 ) ) = '1' else
		0 when ( state_cur(78) and in23 ) = '1' else
		funccall2;
	-- Function 'buf_getb'
	funccall3_next <=
		0 when state_cur(15) = '1' else
		3 when ( state_cur(25) and in6 ) = '1' else
		1 when ( state_cur(30) and in8 ) = '1' else
		2 when state_cur(270) = '1' else
		funccall3;
	-- Function 'buf_getv'
	funccall4_next <=
		0 when state_cur(254) = '1' else
		1 when state_cur(256) = '1' else
		funccall4;
	-- Function 'huff_make_dhuff_tb_ac'
	funccall5_next <=
		0 when state_cur(259) = '1' else
		1 when state_cur(260) = '1' else
		funccall5;
	-- Function 'huff_make_dhuff_tb_dc'
	funccall6_next <=
		1 when state_cur(258) = '1' else
		0 when state_cur(333) = '1' else
		funccall6;
	-- Function 'WriteOneBlock'
	funccall7_next <=
		1 when state_cur(257) = '1' else
		2 when state_cur(445) = '1' else
		3 when state_cur(461) = '1' else
		4 when state_cur(462) = '1' else
		0 when state_cur(469) = '1' else
		funccall7;
	-- Function 'YuvToRgb'
	funccall8_next <=
		0 when state_cur(468) = '1' else
		1 when state_cur(472) = '1' else
		funccall8;
	-- Function 'decode_block'
	funccall9_next <=
		0 when state_cur(418) = '1' else
		1 when state_cur(458) = '1' else
		2 when state_cur(470) = '1' else
		3 when state_cur(471) = '1' else
		funccall9;

	-- Next state bits

	state_next(0) <= (not reset) and ( ( state_cur(422) and in65 ) );
	state_next(1) <= (not reset) and ( state_cur(385) );
	state_next(2) <= (not reset) and ( state_cur(8) or state_cur(3) );
	state_next(3) <= (not reset) and ( ( state_cur(2) and in0 ) );
	state_next(4) <= (not reset) and ( state_cur(377) );
	state_next(5) <= (not reset) and ( ( state_cur(6) and in1 ) );
	state_next(6) <= (not reset) and ( ( state_cur(424) and not ( in67 ) ) );
	state_next(7) <= (not reset) and ( ( state_cur(252) and not ( in49 ) ) or state_cur(202) );
	state_next(8) <= (not reset) and ( ( state_cur(460) and in78 ) or ( state_cur(13) and not ( in2 ) ) or ( state_cur(6) and not ( in1 ) ) );
	state_next(9) <= (not reset) and ( state_cur(327) );
	state_next(10) <= (not reset) and ( state_cur(140) );
	state_next(11) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 16) ) );
	state_next(12) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 15) ) );
	state_next(13) <= (not reset) and ( state_cur(14) or state_cur(7) or state_cur(5) );
	state_next(14) <= (not reset) and ( ( state_cur(17) and not ( in3 ) ) );
	state_next(15) <= (not reset) and ( ( state_cur(13) and in2 ) );
	state_next(16) <= (not reset) and ( ( state_cur(82) and in24 ) );
	state_next(17) <= (not reset) and ( state_cur(19) or state_cur(18) );
	state_next(18) <= (not reset) and ( state_cur(466) or ( state_cur(23) and not ( in4 ) ) );
	state_next(19) <= (not reset) and ( ( state_cur(17) and in3 ) );
	state_next(20) <= (not reset) and ( ( state_cur(454) and in76 ) );
	state_next(21) <= (not reset) and ( ( state_cur(121) and in26 ) );
	state_next(22) <= (not reset) and ( ( state_cur(24) and not ( in5 ) ) );
	state_next(23) <= (not reset) and ( state_cur(159) or state_cur(22) );
	state_next(24) <= (not reset) and ( ( state_cur(25) and not ( in6 ) ) );
	state_next(25) <= (not reset) and ( state_cur(28) or state_cur(26) );
	state_next(26) <= (not reset) and ( ( state_cur(77) and to_stdl(funccall3 = 3) ) or ( state_cur(75) and to_stdl(funccall3 = 3) ) );
	state_next(27) <= (not reset) and ( ( state_cur(29) and not ( in7 ) ) );
	state_next(28) <= (not reset) and ( ( state_cur(77) and to_stdl(funccall3 = 2) ) or ( state_cur(75) and to_stdl(funccall3 = 2) ) );
	state_next(29) <= (not reset) and ( ( state_cur(30) and not ( in8 ) ) );
	state_next(30) <= (not reset) and ( state_cur(32) or state_cur(31) );
	state_next(31) <= (not reset) and ( ( state_cur(77) and to_stdl(funccall3 = 1) ) or ( state_cur(75) and to_stdl(funccall3 = 1) ) );
	state_next(32) <= (not reset) and ( ( state_cur(77) and to_stdl(funccall3 = 0) ) or ( state_cur(75) and to_stdl(funccall3 = 0) ) );
	state_next(33) <= (not reset) and ( state_cur(369) );
	state_next(34) <= (not reset) and ( state_cur(188) or state_cur(38) );
	state_next(35) <= (not reset) and ( ( state_cur(40) and not ( in10 ) ) );
	state_next(36) <= (not reset) and ( state_cur(444) );
	state_next(37) <= (not reset) and ( state_cur(328) );
	state_next(38) <= (not reset) and ( ( state_cur(39) and in9 ) );
	state_next(39) <= (not reset) and ( ( state_cur(40) and in10 ) );
	state_next(40) <= (not reset) and ( state_cur(42) or state_cur(34) );
	state_next(41) <= (not reset) and ( ( state_cur(53) and not ( in14 ) ) );
	state_next(42) <= (not reset) and ( ( state_cur(43) and in11 ) );
	state_next(43) <= (not reset) and ( ( state_cur(427) and not ( in68 ) ) );
	state_next(44) <= (not reset) and ( ( state_cur(45) and not ( in12 ) ) );
	state_next(45) <= (not reset) and ( state_cur(48) or state_cur(46) );
	state_next(46) <= (not reset) and ( ( state_cur(47) and in13 ) );
	state_next(47) <= (not reset) and ( state_cur(49) or state_cur(44) );
	state_next(48) <= (not reset) and ( ( state_cur(45) and in12 ) );
	state_next(49) <= (not reset) and ( ( state_cur(333) ) or ( state_cur(258) ) );
	state_next(50) <= (not reset) and ( state_cur(430) or state_cur(52) );
	state_next(51) <= (not reset) and ( ( state_cur(54) and not ( in15 ) ) );
	state_next(52) <= (not reset) and ( ( state_cur(53) and in14 ) );
	state_next(53) <= (not reset) and ( ( state_cur(54) and in15 ) );
	state_next(54) <= (not reset) and ( state_cur(57) or state_cur(50) );
	state_next(55) <= (not reset) and ( state_cur(372) );
	state_next(56) <= (not reset) and ( state_cur(266) );
	state_next(57) <= (not reset) and ( ( state_cur(59) and in16 ) );
	state_next(58) <= (not reset) and ( state_cur(56) );
	state_next(59) <= (not reset) and ( ( state_cur(366) and not ( in53 ) ) );
	state_next(60) <= (not reset) and ( state_cur(350) );
	state_next(61) <= (not reset) and ( ( state_cur(471) ) or ( state_cur(470) ) or ( state_cur(458) ) or ( state_cur(418) ) );
	state_next(62) <= (not reset) and ( state_cur(208) );
	state_next(63) <= (not reset) and ( ( state_cur(64) and not ( in17 ) ) );
	state_next(64) <= (not reset) and ( state_cur(67) or state_cur(65) );
	state_next(65) <= (not reset) and ( ( state_cur(66) and in18 ) );
	state_next(66) <= (not reset) and ( state_cur(68) or state_cur(63) );
	state_next(67) <= (not reset) and ( ( state_cur(64) and in17 ) );
	state_next(68) <= (not reset) and ( ( state_cur(260) ) or ( state_cur(259) ) );
	state_next(69) <= (not reset) and ( ( state_cur(74) and not ( in21 ) ) );
	state_next(70) <= (not reset) and ( ( state_cur(69) and in19 ) );
	state_next(71) <= (not reset) and ( ( state_cur(80) and to_stdl(funccall2 = 2) ) or ( state_cur(79) and to_stdl(funccall2 = 2) ) );
	state_next(72) <= (not reset) and ( ( state_cur(73) and in20 ) );
	state_next(73) <= (not reset) and ( ( state_cur(74) and in21 ) );
	state_next(74) <= (not reset) and ( state_cur(432) or state_cur(71) );
	state_next(75) <= (not reset) and ( ( state_cur(76) and not ( in22 ) ) );
	state_next(76) <= (not reset) and ( state_cur(81) or ( state_cur(78) and not ( in23 ) ) );
	state_next(77) <= (not reset) and ( ( state_cur(76) and in22 ) );
	state_next(78) <= (not reset) and ( ( state_cur(270) ) or ( state_cur(30) and in8 ) or ( state_cur(25) and in6 ) or ( state_cur(15) ) );
	state_next(79) <= (not reset) and ( ( state_cur(454) and not ( in76 ) ) or ( state_cur(240) and in44 ) );
	state_next(80) <= (not reset) and ( ( state_cur(240) and not ( in44 ) ) );
	state_next(81) <= (not reset) and ( ( state_cur(80) and to_stdl(funccall2 = 0) ) or ( state_cur(79) and to_stdl(funccall2 = 0) ) );
	state_next(82) <= (not reset) and ( state_cur(83) or state_cur(16) );
	state_next(83) <= (not reset) and ( ( state_cur(105) and not ( in25 ) ) );
	state_next(84) <= (not reset) and ( state_cur(302) );
	state_next(85) <= (not reset) and ( state_cur(282) );
	state_next(86) <= (not reset) and ( state_cur(388) );
	state_next(87) <= (not reset) and ( state_cur(122) );
	state_next(88) <= (not reset) and ( state_cur(112) );
	state_next(89) <= (not reset) and ( state_cur(283) );
	state_next(90) <= (not reset) and ( state_cur(89) );
	state_next(91) <= (not reset) and ( state_cur(315) );
	state_next(92) <= (not reset) and ( state_cur(292) );
	state_next(93) <= (not reset) and ( state_cur(99) );
	state_next(94) <= (not reset) and ( state_cur(93) );
	state_next(95) <= (not reset) and ( state_cur(306) );
	state_next(96) <= (not reset) and ( state_cur(317) );
	state_next(97) <= (not reset) and ( state_cur(295) );
	state_next(98) <= (not reset) and ( state_cur(296) );
	state_next(99) <= (not reset) and ( state_cur(290) );
	state_next(100) <= (not reset) and ( state_cur(98) );
	state_next(101) <= (not reset) and ( state_cur(299) );
	state_next(102) <= (not reset) and ( state_cur(106) );
	state_next(103) <= (not reset) and ( state_cur(102) );
	state_next(104) <= (not reset) and ( state_cur(300) );
	state_next(105) <= (not reset) and ( state_cur(224) or state_cur(107) );
	state_next(106) <= (not reset) and ( state_cur(104) );
	state_next(107) <= (not reset) and ( ( state_cur(121) and not ( in26 ) ) );
	state_next(108) <= (not reset) and ( state_cur(307) );
	state_next(109) <= (not reset) and ( state_cur(436) );
	state_next(110) <= (not reset) and ( state_cur(172) );
	state_next(111) <= (not reset) and ( state_cur(314) );
	state_next(112) <= (not reset) and ( state_cur(199) );
	state_next(113) <= (not reset) and ( state_cur(303) );
	state_next(114) <= (not reset) and ( state_cur(111) );
	state_next(115) <= (not reset) and ( state_cur(96) );
	state_next(116) <= (not reset) and ( state_cur(380) );
	state_next(117) <= (not reset) and ( state_cur(345) );
	state_next(118) <= (not reset) and ( state_cur(347) );
	state_next(119) <= (not reset) and ( state_cur(337) );
	state_next(120) <= (not reset) and ( state_cur(180) );
	state_next(121) <= (not reset) and ( state_cur(321) or state_cur(223) );
	state_next(122) <= (not reset) and ( state_cur(183) );
	state_next(123) <= (not reset) and ( ( state_cur(80) and to_stdl(funccall2 = 1) ) or ( state_cur(79) and to_stdl(funccall2 = 1) ) );
	state_next(124) <= (not reset) and ( state_cur(354) );
	state_next(125) <= (not reset) and ( ( state_cur(126) and not ( in32 ) and not ( in31 ) and not ( in30 ) and not ( in29 ) and not ( in28 ) and in27 ) );
	state_next(126) <= (not reset) and ( state_cur(129) or state_cur(128) );
	state_next(127) <= (not reset) and ( state_cur(171) );
	state_next(128) <= (not reset) and ( state_cur(245) );
	state_next(129) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 1) ) );
	state_next(130) <= (not reset) and ( state_cur(234) or ( state_cur(179) and not ( in40 ) ) or ( state_cur(148) and not ( in36 ) ) or state_cur(134) or ( state_cur(126) and not ( in32 ) and not ( in31 ) and not ( in30 ) and not ( in29 ) and not ( in28 ) and not ( in27 ) ) or state_cur(125) );
	state_next(131) <= (not reset) and ( state_cur(273) );
	state_next(132) <= (not reset) and ( ( state_cur(157) and in37 ) );
	state_next(133) <= (not reset) and ( ( state_cur(453) and to_stdl(funccall4 = 0) ) or ( state_cur(131) and to_stdl(funccall4 = 0) ) or ( state_cur(70) and to_stdl(funccall4 = 0) ) );
	state_next(134) <= (not reset) and ( ( state_cur(423) and not ( in66 ) ) );
	state_next(135) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 18) ) );
	state_next(136) <= (not reset) and ( ( state_cur(207) and to_stdl(funccall1 = 6) ) );
	state_next(137) <= (not reset) and ( ( state_cur(138) and in35 ) );
	state_next(138) <= (not reset) and ( state_cur(161) or state_cur(139) );
	state_next(139) <= (not reset) and ( state_cur(136) or state_cur(135) );
	state_next(140) <= (not reset) and ( state_cur(21) );
	state_next(141) <= (not reset) and ( state_cur(331) );
	state_next(142) <= (not reset) and ( state_cur(332) );
	state_next(143) <= (not reset) and ( state_cur(463) );
	state_next(144) <= (not reset) and ( state_cur(9) );
	state_next(145) <= (not reset) and ( state_cur(110) );
	state_next(146) <= (not reset) and ( state_cur(465) );
	state_next(147) <= (not reset) and ( state_cur(10) );
	state_next(148) <= (not reset) and ( state_cur(214) or state_cur(152) );
	state_next(149) <= (not reset) and ( state_cur(319) );
	state_next(150) <= (not reset) and ( state_cur(119) );
	state_next(151) <= (not reset) and ( state_cur(166) );
	state_next(152) <= (not reset) and ( ( state_cur(207) and to_stdl(funccall1 = 5) ) );
	state_next(153) <= (not reset) and ( state_cur(151) );
	state_next(154) <= (not reset) and ( ( state_cur(160) and not ( in38 ) ) );
	state_next(155) <= (not reset) and ( state_cur(341) );
	state_next(156) <= (not reset) and ( state_cur(335) );
	state_next(157) <= (not reset) and ( state_cur(133) );
	state_next(158) <= (not reset) and ( state_cur(186) or ( state_cur(126) and in32 ) );
	state_next(159) <= (not reset) and ( state_cur(167) );
	state_next(160) <= (not reset) and ( state_cur(163) or state_cur(11) );
	state_next(161) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 17) ) );
	state_next(162) <= (not reset) and ( state_cur(156) );
	state_next(163) <= (not reset) and ( ( state_cur(170) and not ( in39 ) ) );
	state_next(164) <= (not reset) and ( ( state_cur(439) and in71 ) );
	state_next(165) <= (not reset) and ( ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 0) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 0) ) );
	state_next(166) <= (not reset) and ( state_cur(361) );
	state_next(167) <= (not reset) and ( ( state_cur(24) and in5 ) );
	state_next(168) <= (not reset) and ( ( state_cur(29) and in7 ) );
	state_next(169) <= (not reset) and ( state_cur(190) or state_cur(187) );
	state_next(170) <= (not reset) and ( state_cur(255) or state_cur(12) );
	state_next(171) <= (not reset) and ( state_cur(87) );
	state_next(172) <= (not reset) and ( state_cur(322) );
	state_next(173) <= (not reset) and ( state_cur(168) );
	state_next(174) <= (not reset) and ( ( state_cur(433) and in70 ) or ( state_cur(59) and not ( in16 ) ) );
	state_next(175) <= (not reset) and ( state_cur(456) );
	state_next(176) <= (not reset) and ( state_cur(348) );
	state_next(177) <= (not reset) and ( state_cur(192) );
	state_next(178) <= (not reset) and ( state_cur(384) );
	state_next(179) <= (not reset) and ( state_cur(184) or state_cur(154) );
	state_next(180) <= (not reset) and ( state_cur(88) );
	state_next(181) <= (not reset) and ( state_cur(455) );
	state_next(182) <= (not reset) and ( state_cur(336) );
	state_next(183) <= (not reset) and ( state_cur(124) );
	state_next(184) <= (not reset) and ( ( state_cur(207) and to_stdl(funccall1 = 4) ) );
	state_next(185) <= (not reset) and ( state_cur(194) );
	state_next(186) <= (not reset) and ( ( state_cur(338) and not ( in52 ) ) );
	state_next(187) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 13) ) );
	state_next(188) <= (not reset) and ( state_cur(426) );
	state_next(189) <= (not reset) and ( state_cur(343) );
	state_next(190) <= (not reset) and ( ( state_cur(212) and not ( in43 ) ) );
	state_next(191) <= (not reset) and ( ( state_cur(252) and in49 ) );
	state_next(192) <= (not reset) and ( state_cur(473) );
	state_next(193) <= (not reset) and ( state_cur(362) );
	state_next(194) <= (not reset) and ( state_cur(176) );
	state_next(195) <= (not reset) and ( state_cur(360) );
	state_next(196) <= (not reset) and ( state_cur(86) );
	state_next(197) <= (not reset) and ( state_cur(55) );
	state_next(198) <= (not reset) and ( state_cur(371) );
	state_next(199) <= (not reset) and ( state_cur(118) );
	state_next(200) <= (not reset) and ( state_cur(376) );
	state_next(201) <= (not reset) and ( state_cur(204) );
	state_next(202) <= (not reset) and ( state_cur(191) );
	state_next(203) <= (not reset) and ( state_cur(359) );
	state_next(204) <= (not reset) and ( state_cur(182) );
	state_next(205) <= (not reset) and ( ( state_cur(210) and not ( in42 ) ) );
	state_next(206) <= (not reset) and ( ( state_cur(210) and in42 ) or ( state_cur(209) and not ( in41 ) ) );
	state_next(207) <= (not reset) and ( state_cur(365) );
	state_next(208) <= (not reset) and ( state_cur(344) );
	state_next(209) <= (not reset) and ( state_cur(213) or state_cur(205) );
	state_next(210) <= (not reset) and ( ( state_cur(209) and in41 ) );
	state_next(211) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 11) ) );
	state_next(212) <= (not reset) and ( state_cur(229) or state_cur(206) );
	state_next(213) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 12) ) );
	state_next(214) <= (not reset) and ( state_cur(353) );
	state_next(215) <= (not reset) and ( state_cur(62) );
	state_next(216) <= (not reset) and ( state_cur(178) );
	state_next(217) <= (not reset) and ( state_cur(389) );
	state_next(218) <= (not reset) and ( state_cur(373) );
	state_next(219) <= (not reset) and ( state_cur(340) );
	state_next(220) <= (not reset) and ( state_cur(374) );
	state_next(221) <= (not reset) and ( state_cur(346) );
	state_next(222) <= (not reset) and ( state_cur(370) );
	state_next(223) <= (not reset) and ( state_cur(367) );
	state_next(224) <= (not reset) and ( state_cur(185) );
	state_next(225) <= (not reset) and ( state_cur(226) );
	state_next(226) <= (not reset) and ( state_cur(227) );
	state_next(227) <= (not reset) and ( state_cur(218) );
	state_next(228) <= (not reset) and ( state_cur(230) );
	state_next(229) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 10) ) );
	state_next(230) <= (not reset) and ( state_cur(225) );
	state_next(231) <= (not reset) and ( state_cur(233) );
	state_next(232) <= (not reset) and ( state_cur(280) );
	state_next(233) <= (not reset) and ( state_cur(232) );
	state_next(234) <= (not reset) and ( ( state_cur(241) and not ( in45 ) ) );
	state_next(235) <= (not reset) and ( state_cur(164) );
	state_next(236) <= (not reset) and ( state_cur(165) );
	state_next(237) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 8) ) );
	state_next(238) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 7) ) );
	state_next(239) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 9) ) );
	state_next(240) <= (not reset) and ( state_cur(20) );
	state_next(241) <= (not reset) and ( state_cur(247) or state_cur(239) );
	state_next(242) <= (not reset) and ( ( state_cur(241) and in45 ) );
	state_next(243) <= (not reset) and ( ( state_cur(207) and to_stdl(funccall1 = 2) ) );
	state_next(244) <= (not reset) and ( ( state_cur(207) and to_stdl(funccall1 = 1) ) );
	state_next(245) <= (not reset) and ( ( state_cur(246) and in46 ) );
	state_next(246) <= (not reset) and ( ( state_cur(251) and not ( in48 ) ) );
	state_next(247) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 6) ) );
	state_next(248) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 3) ) );
	state_next(249) <= (not reset) and ( state_cur(250) or state_cur(248) );
	state_next(250) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 2) ) );
	state_next(251) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 4) ) );
	state_next(252) <= (not reset) and ( state_cur(253) );
	state_next(253) <= (not reset) and ( ( state_cur(453) and to_stdl(funccall4 = 1) ) or ( state_cur(131) and to_stdl(funccall4 = 1) ) or ( state_cur(70) and to_stdl(funccall4 = 1) ) );
	state_next(254) <= (not reset) and ( ( state_cur(23) and in4 ) );
	state_next(255) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 14) ) );
	state_next(256) <= (not reset) and ( ( state_cur(460) and not ( in78 ) ) );
	state_next(257) <= (not reset) and ( ( state_cur(399) and in56 ) );
	state_next(258) <= (not reset) and ( ( state_cur(35) and to_stdl(funccall6 = 0) ) );
	state_next(259) <= (not reset) and ( ( state_cur(35) and to_stdl(funccall6 = 1) ) );
	state_next(260) <= (not reset) and ( ( state_cur(51) and to_stdl(funccall5 = 0) ) );
	state_next(261) <= (not reset) and ( ( state_cur(51) and to_stdl(funccall5 = 1) ) );
	state_next(262) <= (not reset) and ( state_cur(391) or ( state_cur(262) and not (in50) ) );
	state_next(263) <= (not reset) and ( ( state_cur(392) and not ( in55 ) ) or ( state_cur(263) and not (in50) ) );
	state_next(264) <= (not reset) and ( state_cur(386) or ( state_cur(264) and not (in50) ) );
	state_next(265) <= (not reset) and ( ( state_cur(423) and in66 ) or state_cur(397) or ( state_cur(265) and not (in51) ) );
	state_next(266) <= (not reset) and ( state_cur(85) );
	state_next(267) <= (not reset) and ( state_cur(58) );
	state_next(268) <= (not reset) and ( state_cur(267) );
	state_next(269) <= (not reset) and ( state_cur(268) );
	state_next(270) <= (not reset) and ( state_cur(61) );
	state_next(271) <= (not reset) and ( ( state_cur(256) ) or ( state_cur(254) ) );
	state_next(272) <= (not reset) and ( state_cur(198) );
	state_next(273) <= (not reset) and ( ( state_cur(69) and not ( in19 ) ) );
	state_next(274) <= (not reset) and ( state_cur(272) );
	state_next(275) <= (not reset) and ( ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 4) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 4) ) );
	state_next(276) <= (not reset) and ( state_cur(275) );
	state_next(277) <= (not reset) and ( state_cur(269) );
	state_next(278) <= (not reset) and ( state_cur(277) );
	state_next(279) <= (not reset) and ( state_cur(274) );
	state_next(280) <= (not reset) and ( state_cur(279) );
	state_next(281) <= (not reset) and ( state_cur(84) );
	state_next(282) <= (not reset) and ( state_cur(281) );
	state_next(283) <= (not reset) and ( state_cur(92) );
	state_next(284) <= (not reset) and ( state_cur(90) );
	state_next(285) <= (not reset) and ( state_cur(284) );
	state_next(286) <= (not reset) and ( state_cur(285) );
	state_next(287) <= (not reset) and ( state_cur(286) );
	state_next(288) <= (not reset) and ( state_cur(287) );
	state_next(289) <= (not reset) and ( state_cur(288) );
	state_next(290) <= (not reset) and ( state_cur(289) );
	state_next(291) <= (not reset) and ( state_cur(91) );
	state_next(292) <= (not reset) and ( state_cur(291) );
	state_next(293) <= (not reset) and ( state_cur(94) );
	state_next(294) <= (not reset) and ( state_cur(293) );
	state_next(295) <= (not reset) and ( state_cur(294) );
	state_next(296) <= (not reset) and ( state_cur(97) );
	state_next(297) <= (not reset) and ( state_cur(100) );
	state_next(298) <= (not reset) and ( state_cur(297) );
	state_next(299) <= (not reset) and ( state_cur(298) );
	state_next(300) <= (not reset) and ( state_cur(101) );
	state_next(301) <= (not reset) and ( state_cur(103) );
	state_next(302) <= (not reset) and ( state_cur(301) );
	state_next(303) <= (not reset) and ( state_cur(357) );
	state_next(304) <= (not reset) and ( state_cur(434) );
	state_next(305) <= (not reset) and ( state_cur(425) );
	state_next(306) <= (not reset) and ( state_cur(305) );
	state_next(307) <= (not reset) and ( state_cur(304) );
	state_next(308) <= (not reset) and ( state_cur(108) );
	state_next(309) <= (not reset) and ( state_cur(308) );
	state_next(310) <= (not reset) and ( state_cur(95) );
	state_next(311) <= (not reset) and ( state_cur(310) );
	state_next(312) <= (not reset) and ( state_cur(311) );
	state_next(313) <= (not reset) and ( state_cur(309) );
	state_next(314) <= (not reset) and ( state_cur(313) );
	state_next(315) <= (not reset) and ( state_cur(114) );
	state_next(316) <= (not reset) and ( state_cur(318) );
	state_next(317) <= (not reset) and ( state_cur(312) );
	state_next(318) <= (not reset) and ( state_cur(329) );
	state_next(319) <= (not reset) and ( state_cur(316) );
	state_next(320) <= (not reset) and ( state_cur(326) );
	state_next(321) <= (not reset) and ( state_cur(115) );
	state_next(322) <= (not reset) and ( state_cur(320) );
	state_next(323) <= (not reset) and ( state_cur(330) );
	state_next(324) <= (not reset) and ( ( state_cur(78) and in23 ) or ( state_cur(73) and not ( in20 ) ) or ( state_cur(72) ) );
	state_next(325) <= (not reset) and ( state_cur(323) );
	state_next(326) <= (not reset) and ( state_cur(325) );
	state_next(327) <= (not reset) and ( state_cur(155) );
	state_next(328) <= (not reset) and ( state_cur(145) );
	state_next(329) <= (not reset) and ( state_cur(141) );
	state_next(330) <= (not reset) and ( state_cur(142) );
	state_next(331) <= (not reset) and ( state_cur(113) );
	state_next(332) <= (not reset) and ( state_cur(438) );
	state_next(333) <= (not reset) and ( state_cur(158) );
	state_next(334) <= (not reset) and ( state_cur(197) );
	state_next(335) <= (not reset) and ( state_cur(189) );
	state_next(336) <= (not reset) and ( state_cur(203) );
	state_next(337) <= (not reset) and ( state_cur(358) );
	state_next(338) <= (not reset) and ( state_cur(169) );
	state_next(339) <= (not reset) and ( state_cur(349) );
	state_next(340) <= (not reset) and ( state_cur(177) );
	state_next(341) <= (not reset) and ( state_cur(339) );
	state_next(342) <= (not reset) and ( state_cur(382) );
	state_next(343) <= (not reset) and ( state_cur(150) );
	state_next(344) <= (not reset) and ( state_cur(442) );
	state_next(345) <= (not reset) and ( state_cur(400) );
	state_next(346) <= (not reset) and ( state_cur(200) );
	state_next(347) <= (not reset) and ( state_cur(162) );
	state_next(348) <= (not reset) and ( state_cur(193) );
	state_next(349) <= (not reset) and ( state_cur(219) );
	state_next(350) <= (not reset) and ( state_cur(37) );
	state_next(351) <= (not reset) and ( state_cur(404) );
	state_next(352) <= (not reset) and ( state_cur(1) );
	state_next(353) <= (not reset) and ( ( state_cur(138) and not ( in35 ) ) );
	state_next(354) <= (not reset) and ( ( state_cur(105) and in25 ) );
	state_next(355) <= (not reset) and ( state_cur(175) );
	state_next(356) <= (not reset) and ( state_cur(4) );
	state_next(357) <= (not reset) and ( ( state_cur(82) and not ( in24 ) ) );
	state_next(358) <= (not reset) and ( state_cur(117) );
	state_next(359) <= (not reset) and ( state_cur(352) );
	state_next(360) <= (not reset) and ( state_cur(368) );
	state_next(361) <= (not reset) and ( state_cur(33) );
	state_next(362) <= (not reset) and ( state_cur(356) );
	state_next(363) <= (not reset) and ( ( state_cur(451) and in74 ) );
	state_next(364) <= (not reset) and ( state_cur(228) );
	state_next(365) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 5) ) or ( state_cur(244) ) or ( state_cur(137) and in34 ) or ( state_cur(126) and not ( in32 ) and not ( in31 ) and not ( in30 ) and not ( in29 ) and in28 ) or ( state_cur(126) and not ( in32 ) and not ( in31 ) and not ( in30 ) and in29 ) or ( state_cur(126) and not ( in32 ) and not ( in31 ) and in30 ) or ( state_cur(126) and not ( in32 ) and in31 ) );
	state_next(366) <= (not reset) and ( state_cur(441) );
	state_next(367) <= (not reset) and ( state_cur(201) );
	state_next(368) <= (not reset) and ( state_cur(221) );
	state_next(369) <= (not reset) and ( state_cur(231) );
	state_next(370) <= (not reset) and ( state_cur(394) );
	state_next(371) <= (not reset) and ( ( state_cur(2) and not ( in0 ) ) );
	state_next(372) <= (not reset) and ( state_cur(375) );
	state_next(373) <= (not reset) and ( state_cur(215) );
	state_next(374) <= (not reset) and ( state_cur(217) );
	state_next(375) <= (not reset) and ( state_cur(355) );
	state_next(376) <= (not reset) and ( state_cur(381) );
	state_next(377) <= (not reset) and ( state_cur(127) );
	state_next(378) <= (not reset) and ( ( state_cur(428) and in69 ) or ( state_cur(43) and not ( in11 ) ) );
	state_next(379) <= (not reset) and ( ( state_cur(47) and not ( in13 ) ) );
	state_next(380) <= (not reset) and ( state_cur(351) );
	state_next(381) <= (not reset) and ( state_cur(216) );
	state_next(382) <= (not reset) and ( state_cur(195) );
	state_next(383) <= (not reset) and ( ( state_cur(469) ) or ( state_cur(462) ) or ( state_cur(461) ) or ( state_cur(445) ) or ( state_cur(257) ) );
	state_next(384) <= (not reset) and ( state_cur(196) );
	state_next(385) <= (not reset) and ( state_cur(120) );
	state_next(386) <= (not reset) and ( ( state_cur(263) and not ( not (in50) ) ) );
	state_next(387) <= (not reset) and ( state_cur(342) );
	state_next(388) <= (not reset) and ( state_cur(60) );
	state_next(389) <= (not reset) and ( state_cur(235) );
	state_next(390) <= (not reset) and ( ( state_cur(262) and not ( not (in50) ) ) );
	state_next(391) <= (not reset) and ( state_cur(393) or ( state_cur(390) and in54 ) );
	state_next(392) <= (not reset) and ( ( state_cur(390) and not ( in54 ) ) );
	state_next(393) <= (not reset) and ( state_cur(395) or ( state_cur(392) and in55 ) );
	state_next(394) <= (not reset) and ( state_cur(364) );
	state_next(395) <= (not reset) and ( ( state_cur(416) and not ( in62 ) ) or ( state_cur(409) and not ( in59 ) ) );
	state_next(396) <= (not reset) and ( ( state_cur(396) and to_stdl(funccall0 = 0) ) or ( state_cur(338) and in52 ) or ( state_cur(251) and in48 ) or ( state_cur(249) and not ( in47 ) ) or ( state_cur(249) and in47 ) or ( state_cur(246) and not ( in46 ) ) or ( state_cur(243) ) or ( state_cur(242) ) or ( state_cur(238) ) or ( state_cur(237) ) or ( state_cur(212) and in43 ) or ( state_cur(211) ) or ( state_cur(207) and to_stdl(funccall1 = 0) ) or ( state_cur(207) and to_stdl(funccall1 = 3) ) or ( state_cur(179) and in40 ) or ( state_cur(170) and in39 ) or ( state_cur(160) and in38 ) or ( state_cur(148) and in36 ) or ( state_cur(137) and not ( in34 ) ) or ( state_cur(130) and not ( in33 ) ) or ( state_cur(130) and in33 ) );
	state_next(397) <= (not reset) and ( ( state_cur(457) and not ( not (in77) ) ) or ( state_cur(264) and not ( not (in50) ) ) );
	state_next(398) <= (not reset) and ( ( state_cur(399) and not ( in56 ) ) );
	state_next(399) <= (not reset) and ( state_cur(401) or state_cur(276) );
	state_next(400) <= (not reset) and ( state_cur(109) );
	state_next(401) <= (not reset) and ( ( state_cur(403) and not ( in57 ) ) );
	state_next(402) <= (not reset) and ( ( state_cur(439) and not ( in71 ) and to_stdl(funccall8 = 1) ) );
	state_next(403) <= (not reset) and ( state_cur(405) or state_cur(402) );
	state_next(404) <= (not reset) and ( state_cur(387) );
	state_next(405) <= (not reset) and ( ( state_cur(278) and to_stdl(funccall9 = 3) ) );
	state_next(406) <= (not reset) and ( ( state_cur(278) and to_stdl(funccall9 = 1) ) );
	state_next(407) <= (not reset) and ( state_cur(408) or state_cur(406) );
	state_next(408) <= (not reset) and ( ( state_cur(409) and in59 ) );
	state_next(409) <= (not reset) and ( ( state_cur(417) and not ( in63 ) ) or state_cur(398) );
	state_next(410) <= (not reset) and ( ( state_cur(411) and not ( in60 ) ) );
	state_next(411) <= (not reset) and ( state_cur(412) or state_cur(236) );
	state_next(412) <= (not reset) and ( ( state_cur(439) and not ( in71 ) and to_stdl(funccall8 = 0) ) );
	state_next(413) <= (not reset) and ( ( state_cur(278) and to_stdl(funccall9 = 0) ) );
	state_next(414) <= (not reset) and ( state_cur(415) or state_cur(413) );
	state_next(415) <= (not reset) and ( ( state_cur(416) and in62 ) );
	state_next(416) <= (not reset) and ( ( state_cur(417) and in63 ) or state_cur(410) );
	state_next(417) <= (not reset) and ( ( state_cur(419) and not ( in64 ) ) );
	state_next(418) <= (not reset) and ( ( state_cur(414) and in61 ) );
	state_next(419) <= (not reset) and ( state_cur(421) or state_cur(420) );
	state_next(420) <= (not reset) and ( ( state_cur(419) and in64 ) );
	state_next(421) <= (not reset) and ( ( state_cur(422) and not ( in65 ) ) );
	state_next(422) <= (not reset) and ( state_cur(261) or state_cur(0) );
	state_next(423) <= (not reset) and ( ( state_cur(265) and not ( not (in51) ) ) );
	state_next(424) <= (not reset) and ( state_cur(435) );
	state_next(425) <= (not reset) and ( state_cur(146) );
	state_next(426) <= (not reset) and ( ( state_cur(39) and not ( in9 ) ) );
	state_next(427) <= (not reset) and ( state_cur(429) );
	state_next(428) <= (not reset) and ( state_cur(378) );
	state_next(429) <= (not reset) and ( state_cur(431) or ( state_cur(428) and not ( in69 ) ) or ( state_cur(427) and in68 ) );
	state_next(430) <= (not reset) and ( state_cur(41) );
	state_next(431) <= (not reset) and ( state_cur(379) );
	state_next(432) <= (not reset) and ( state_cur(271) );
	state_next(433) <= (not reset) and ( state_cur(174) );
	state_next(434) <= (not reset) and ( state_cur(143) );
	state_next(435) <= (not reset) and ( state_cur(173) or state_cur(27) );
	state_next(436) <= (not reset) and ( state_cur(181) );
	state_next(437) <= (not reset) and ( state_cur(443) or ( state_cur(157) and not ( in37 ) ) );
	state_next(438) <= (not reset) and ( state_cur(334) );
	state_next(439) <= (not reset) and ( state_cur(440) or state_cur(220) );
	state_next(440) <= (not reset) and ( ( state_cur(472) ) or ( state_cur(468) ) );
	state_next(441) <= (not reset) and ( ( state_cur(433) and not ( in70 ) ) or ( state_cur(366) and in53 ) or state_cur(36) );
	state_next(442) <= (not reset) and ( state_cur(153) );
	state_next(443) <= (not reset) and ( state_cur(132) );
	state_next(444) <= (not reset) and ( ( state_cur(66) and not ( in18 ) ) );
	state_next(445) <= (not reset) and ( ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 1) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 1) ) );
	state_next(446) <= (not reset) and ( ( state_cur(449) and not ( in73 ) ) or ( state_cur(448) and not ( in72 ) ) );
	state_next(447) <= (not reset) and ( state_cur(450) );
	state_next(448) <= (not reset) and ( ( state_cur(449) and in73 ) );
	state_next(449) <= (not reset) and ( state_cur(447) or state_cur(363) );
	state_next(450) <= (not reset) and ( ( state_cur(448) and in72 ) );
	state_next(451) <= (not reset) and ( ( state_cur(452) and in75 ) );
	state_next(452) <= (not reset) and ( state_cur(446) or state_cur(383) );
	state_next(453) <= (not reset) and ( state_cur(123) );
	state_next(454) <= (not reset) and ( state_cur(324) );
	state_next(455) <= (not reset) and ( state_cur(222) );
	state_next(456) <= (not reset) and ( state_cur(149) );
	state_next(457) <= reset or ( ( state_cur(457) and not (in77) ) );
	state_next(458) <= (not reset) and ( ( state_cur(407) and in58 ) );
	state_next(459) <= (not reset) and ( ( state_cur(424) and in67 ) );
	state_next(460) <= (not reset) and ( state_cur(459) );
	state_next(461) <= (not reset) and ( ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 2) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 2) ) );
	state_next(462) <= (not reset) and ( ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 3) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 3) ) );
	state_next(463) <= (not reset) and ( state_cur(464) );
	state_next(464) <= (not reset) and ( state_cur(144) );
	state_next(465) <= (not reset) and ( state_cur(467) );
	state_next(466) <= (not reset) and ( state_cur(437) );
	state_next(467) <= (not reset) and ( state_cur(147) );
	state_next(468) <= (not reset) and ( ( state_cur(414) and not ( in61 ) ) );
	state_next(469) <= (not reset) and ( ( state_cur(411) and in60 ) );
	state_next(470) <= (not reset) and ( ( state_cur(407) and not ( in58 ) ) );
	state_next(471) <= (not reset) and ( ( state_cur(278) and to_stdl(funccall9 = 2) ) );
	state_next(472) <= (not reset) and ( ( state_cur(403) and in57 ) );
	state_next(473) <= (not reset) and ( state_cur(116) );

	-- Assignment of buffers for buffered outputs

	out1057_bufn <= state_cur(127) or state_cur(425);
	out59_bufn <= state_cur(305) or state_cur(377);
	out447_bufn <= state_cur(382) or state_cur(111);
	out157_bufn <= state_cur(28) or state_cur(26) or ( state_cur(25) and not ( in6 ) );
	out450_bufn <= state_cur(194) or state_cur(96);
	out1012_bufn <= state_cur(221) or state_cur(291);
	out1072_bufn <= state_cur(351) or state_cur(308);
	out999_bufn <= state_cur(196) or state_cur(286);
	out437_bufn <= state_cur(94) or state_cur(172);
	out415_bufn <= state_cur(330) or state_cur(98);
	out426_bufn <= state_cur(321) or state_cur(223) or state_cur(224) or state_cur(107);
	out375_bufn <= state_cur(360) or state_cur(315);
	out704_bufn <= state_cur(356) or state_cur(193) or state_cur(311) or state_cur(310) or state_cur(95) or state_cur(362);
	out973_bufn <= state_cur(275) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 4) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 4) );
	out11_bufn <= state_cur(222) or state_cur(153) or state_cur(181) or state_cur(109) or state_cur(364) or state_cur(120) or state_cur(215) or state_cur(394) or state_cur(231) or state_cur(201) or state_cur(228) or state_cur(33) or state_cur(352) or state_cur(117) or state_cur(1) or state_cur(162) or state_cur(400) or state_cur(442) or state_cur(150) or state_cur(358) or state_cur(203) or state_cur(189) or state_cur(279) or state_cur(274) or state_cur(272) or state_cur(198) or state_cur(232) or state_cur(280) or state_cur(233) or state_cur(225) or state_cur(230) or state_cur(218) or state_cur(227) or state_cur(226) or state_cur(367) or state_cur(370) or state_cur(373) or state_cur(62) or state_cur(344) or state_cur(182) or state_cur(359) or state_cur(204) or state_cur(118) or state_cur(371) or state_cur(343) or state_cur(336) or state_cur(455) or state_cur(88) or state_cur(361) or state_cur(156) or state_cur(335) or state_cur(151) or state_cur(166) or state_cur(119) or state_cur(180) or state_cur(337) or state_cur(347) or state_cur(345) or state_cur(199) or state_cur(436) or state_cur(112) or state_cur(208) or state_cur(369) or state_cur(385);
	out549_bufn <= state_cur(87) or state_cur(465);
	out453_bufn <= state_cur(304) or state_cur(380);
	out1231_bufn <= state_cur(261) or state_cur(0) or state_cur(421) or state_cur(420) or state_cur(415) or state_cur(413) or state_cur(412) or state_cur(236) or state_cur(408) or state_cur(406) or state_cur(405) or state_cur(402) or state_cur(401) or state_cur(276);
	out87_bufn <= state_cur(147) or state_cur(467) or state_cur(312) or state_cur(10) or state_cur(465) or state_cur(21) or state_cur(96) or state_cur(317) or state_cur(140);
	out401_bufn <= state_cur(4) or state_cur(306);
	out990_bufn <= state_cur(316) or state_cur(281);
	out378_bufn <= state_cur(376) or state_cur(292);
	out1302_bufn <= state_cur(132) or state_cur(443) or ( state_cur(157) and not ( in37 ) );
	out27_bufn <= ( state_cur(448) and in72 ) or ( state_cur(433) and not ( in70 ) ) or ( state_cur(366) and in53 ) or state_cur(36) or state_cur(431) or ( state_cur(428) and not ( in69 ) ) or ( state_cur(427) and in68 ) or state_cur(193) or state_cur(311) or state_cur(310) or state_cur(95) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 4) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 4) ) or state_cur(362) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 0) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 0) ) or state_cur(186) or ( state_cur(126) and in32 ) or state_cur(136) or state_cur(135) or ( state_cur(64) and in17 ) or ( state_cur(45) and in12 ) or ( state_cur(77) and to_stdl(funccall3 = 1) ) or ( state_cur(75) and to_stdl(funccall3 = 1) ) or ( state_cur(77) and to_stdl(funccall3 = 3) ) or ( state_cur(75) and to_stdl(funccall3 = 3) ) or ( state_cur(2) and in0 );
	out569_bufn <= ( state_cur(138) and not ( in35 ) ) or ( state_cur(207) and to_stdl(funccall1 = 5) );
	out1030_bufn <= state_cur(438) or state_cur(101);
	out537_bufn <= state_cur(293) or state_cur(110);
	out77_bufn <= state_cur(144) or state_cur(464) or state_cur(143) or state_cur(155) or state_cur(114) or state_cur(313) or state_cur(309) or state_cur(308) or state_cur(108) or state_cur(304) or state_cur(434) or state_cur(301) or state_cur(103) or state_cur(101) or state_cur(298) or state_cur(297) or state_cur(100) or state_cur(97) or state_cur(294) or state_cur(293) or state_cur(94) or state_cur(291) or state_cur(91) or state_cur(289) or state_cur(288) or state_cur(287) or state_cur(286) or state_cur(285) or state_cur(284) or state_cur(90) or state_cur(92) or state_cur(281) or state_cur(84) or state_cur(277) or state_cur(269) or state_cur(268) or state_cur(267) or state_cur(58) or state_cur(85) or state_cur(9) or state_cur(463) or state_cur(111) or state_cur(314) or state_cur(307) or state_cur(104) or state_cur(300) or state_cur(102) or state_cur(106) or state_cur(299) or state_cur(98) or state_cur(290) or state_cur(296) or state_cur(295) or state_cur(93) or state_cur(99) or state_cur(292) or state_cur(315) or state_cur(89) or state_cur(283) or state_cur(282) or state_cur(302) or state_cur(56) or state_cur(266) or state_cur(327);
	out1318_bufn <= ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 3) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 3) ) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 1) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 1) );
	out533_bufn <= state_cur(219) or state_cur(9);
	out32_bufn <= state_cur(305) or state_cur(176) or state_cur(317) or state_cur(377);
	out1027_bufn <= state_cur(142) or state_cur(298);
	out599_bufn <= ( state_cur(35) and to_stdl(funccall6 = 0) ) or state_cur(186) or ( state_cur(126) and in32 );
	out668_bufn <= state_cur(84) or state_cur(456);
	out568_bufn <= state_cur(261) or state_cur(0) or state_cur(421) or state_cur(420) or state_cur(415) or state_cur(413) or state_cur(412) or state_cur(236) or state_cur(401) or state_cur(276) or ( state_cur(207) and to_stdl(funccall1 = 4) ) or ( state_cur(207) and to_stdl(funccall1 = 5) );
	out225_bufn <= ( state_cur(39) and not ( in9 ) ) or ( state_cur(53) and not ( in14 ) );
	out700_bufn <= state_cur(143) or state_cur(473);
	out638_bufn <= ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 4) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 4) ) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 0) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 0) );
	out670_bufn <= state_cur(312) or state_cur(348);
	out433_bufn <= state_cur(116) or state_cur(307);
	out896_bufn <= ( state_cur(411) and in60 ) or ( state_cur(399) and in56 );
	out575_bufn <= state_cur(163) or state_cur(11) or ( state_cur(160) and not ( in38 ) );
	out428_bufn <= state_cur(197) or state_cur(104);
	out72_bufn <= state_cur(144) or state_cur(464) or state_cur(143) or state_cur(155) or state_cur(114) or state_cur(313) or state_cur(309) or state_cur(308) or state_cur(108) or state_cur(304) or state_cur(434) or state_cur(301) or state_cur(103) or state_cur(101) or state_cur(298) or state_cur(297) or state_cur(100) or state_cur(97) or state_cur(294) or state_cur(293) or state_cur(94) or state_cur(291) or state_cur(91) or state_cur(289) or state_cur(288) or state_cur(287) or state_cur(286) or state_cur(285) or state_cur(284) or state_cur(90) or state_cur(92) or state_cur(281) or state_cur(84) or state_cur(277) or state_cur(269) or state_cur(268) or state_cur(267) or state_cur(58) or state_cur(85) or state_cur(9) or state_cur(463) or state_cur(111) or state_cur(314) or state_cur(307) or state_cur(104) or state_cur(300) or state_cur(102) or state_cur(106) or state_cur(299) or state_cur(98) or state_cur(290) or state_cur(296) or state_cur(295) or state_cur(93) or state_cur(99) or state_cur(292) or state_cur(315) or state_cur(89) or state_cur(283) or state_cur(282) or state_cur(302) or state_cur(56) or state_cur(266) or ( state_cur(82) and in24 ) or state_cur(327);
	out404_bufn <= state_cur(115) or state_cur(312) or state_cur(185) or state_cur(176) or state_cur(194) or state_cur(348) or state_cur(96) or state_cur(317);
	out98_bufn <= ( state_cur(396) and to_stdl(funccall0 = 15) ) or ( state_cur(396) and to_stdl(funccall0 = 16) );
	out67_bufn <= ( state_cur(424) and in67 ) or ( state_cur(252) and not ( in49 ) ) or state_cur(202);
	out635_bufn <= state_cur(165) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 0) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 0) );
	out381_bufn <= state_cur(145) or state_cur(99);
	out222_bufn <= ( state_cur(433) and not ( in70 ) ) or ( state_cur(366) and in53 ) or state_cur(36) or state_cur(41) or ( state_cur(64) and in17 ) or ( state_cur(53) and not ( in14 ) );
	out339_bufn <= state_cur(273) or ( state_cur(76) and in22 ) or ( state_cur(76) and not ( in22 ) );
	out268_bufn <= state_cur(41) or ( state_cur(53) and in14 );
	out419_bufn <= state_cur(375) or state_cur(106);
	out559_bufn <= ( state_cur(138) and not ( in35 ) ) or state_cur(353) or state_cur(214) or state_cur(152);
	out1002_bufn <= state_cur(60) or state_cur(287);
	out1006_bufn <= state_cur(37) or state_cur(289);
	out276_bufn <= state_cur(318) or state_cur(266);
	out205_bufn <= state_cur(116) or state_cur(149) or state_cur(334) or state_cur(387) or state_cur(60) or state_cur(342) or state_cur(196) or state_cur(195) or state_cur(216) or state_cur(351) or state_cur(381) or state_cur(355) or state_cur(375) or state_cur(221) or state_cur(368) or ( state_cur(82) and not ( in24 ) ) or state_cur(175) or state_cur(404) or state_cur(37) or state_cur(219) or state_cur(200) or state_cur(382) or state_cur(339) or state_cur(177) or state_cur(349) or state_cur(197) or state_cur(438) or state_cur(113) or state_cur(142) or state_cur(141) or state_cur(145) or state_cur(325) or state_cur(323) or state_cur(330) or state_cur(320) or state_cur(326) or state_cur(316) or state_cur(329) or state_cur(318) or state_cur(357) or state_cur(346) or state_cur(340) or state_cur(178) or state_cur(376) or state_cur(55) or state_cur(86) or state_cur(360) or state_cur(473) or state_cur(384) or state_cur(192) or state_cur(456) or state_cur(322) or state_cur(341) or state_cur(319) or state_cur(110) or state_cur(332) or state_cur(331) or state_cur(380) or state_cur(303) or state_cur(172) or state_cur(388) or state_cur(350) or state_cur(372) or state_cur(328);
	out943_bufn <= state_cur(329) or state_cur(85);
	out1080_bufn <= state_cur(193) or state_cur(311);
	out408_bufn <= state_cur(322) or state_cur(295);
	out252_bufn <= state_cur(431) or ( state_cur(428) and not ( in69 ) ) or ( state_cur(427) and in68 ) or ( state_cur(39) and not ( in9 ) ) or state_cur(426) or ( state_cur(45) and in12 );
	out71_bufn <= state_cur(341) or state_cur(327);
	out672_bufn <= state_cur(434) or state_cur(192);
	out357_bufn <= state_cur(319) or state_cur(282);
	out441_bufn <= state_cur(195) or state_cur(314);
	out1084_bufn <= state_cur(387) or state_cur(313);
	out144_bufn <= ( state_cur(78) and in23 ) or ( state_cur(73) and not ( in20 ) ) or ( state_cur(72) ) or ( state_cur(454) and in76 );
	out574_bufn <= state_cur(184) or state_cur(154) or ( state_cur(170) and not ( in39 ) ) or ( state_cur(160) and not ( in38 ) );
	out210_bufn <= ( state_cur(39) and not ( in9 ) ) or ( state_cur(40) and in10 );
	out128_bufn <= state_cur(306) or ( state_cur(82) and in24 );
	out360_bufn <= state_cur(288) or state_cur(388);
	out948_bufn <= state_cur(141) or state_cur(58);
	out506_bufn <= ( state_cur(453) and to_stdl(funccall4 = 1) ) or ( state_cur(131) and to_stdl(funccall4 = 1) ) or ( state_cur(70) and to_stdl(funccall4 = 1) ) or ( state_cur(453) and to_stdl(funccall4 = 0) ) or ( state_cur(131) and to_stdl(funccall4 = 0) ) or ( state_cur(70) and to_stdl(funccall4 = 0) );
	out207_bufn <= state_cur(93) or state_cur(328);
	out1083_bufn <= state_cur(342) or state_cur(309);
	out491_bufn <= state_cur(146) or state_cur(171);
	out4_bufn <= state_cur(147) or state_cur(467) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 3) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 3) ) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 2) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 2) ) or state_cur(446) or state_cur(383) or state_cur(447) or state_cur(363) or state_cur(450) or ( state_cur(449) and not ( in73 ) ) or ( state_cur(448) and not ( in72 ) ) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 1) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 1) ) or state_cur(132) or ( state_cur(433) and not ( in70 ) ) or ( state_cur(366) and in53 ) or state_cur(36) or state_cur(41) or state_cur(431) or ( state_cur(428) and not ( in69 ) ) or ( state_cur(427) and in68 ) or state_cur(146) or ( state_cur(265) and not ( not (in51) ) ) or ( state_cur(419) and in64 ) or ( state_cur(278) and to_stdl(funccall9 = 0) ) or ( state_cur(411) and not ( in60 ) ) or ( state_cur(278) and to_stdl(funccall9 = 1) ) or ( state_cur(439) and not ( in71 ) and to_stdl(funccall8 = 1) ) or ( state_cur(399) and not ( in56 ) ) or ( state_cur(396) and to_stdl(funccall0 = 0) ) or ( state_cur(338) and in52 ) or ( state_cur(251) and in48 ) or ( state_cur(249) and not ( in47 ) ) or ( state_cur(249) and in47 ) or ( state_cur(246) and not ( in46 ) ) or ( state_cur(243) ) or ( state_cur(242) ) or ( state_cur(238) ) or ( state_cur(237) ) or ( state_cur(212) and in43 ) or ( state_cur(211) ) or ( state_cur(207) and to_stdl(funccall1 = 0) ) or ( state_cur(207) and to_stdl(funccall1 = 3) ) or ( state_cur(179) and in40 ) or ( state_cur(170) and in39 ) or ( state_cur(160) and in38 ) or ( state_cur(148) and in36 ) or ( state_cur(137) and not ( in34 ) ) or ( state_cur(130) and not ( in33 ) ) or ( state_cur(130) and in33 ) or ( state_cur(390) and not ( in54 ) ) or ( state_cur(262) and not ( not (in50) ) ) or ( state_cur(428) and in69 ) or ( state_cur(43) and not ( in11 ) ) or ( state_cur(2) and not ( in0 ) ) or ( state_cur(396) and to_stdl(funccall0 = 5) ) or ( state_cur(244) ) or ( state_cur(137) and in34 ) or ( state_cur(126) and not ( in32 ) and not ( in31 ) and not ( in30 ) and not ( in29 ) and in28 ) or ( state_cur(126) and not ( in32 ) and not ( in31 ) and not ( in30 ) and in29 ) or ( state_cur(126) and not ( in32 ) and not ( in31 ) and in30 ) or ( state_cur(126) and not ( in32 ) and in31 ) or ( state_cur(105) and in25 ) or ( state_cur(78) and in23 ) or ( state_cur(73) and not ( in20 ) ) or ( state_cur(72) ) or state_cur(312) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 4) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 4) ) or ( state_cur(396) and to_stdl(funccall0 = 9) ) or state_cur(164) or state_cur(374) or state_cur(365) or ( state_cur(210) and in42 ) or ( state_cur(209) and not ( in41 ) ) or ( state_cur(210) and not ( in42 ) ) or state_cur(191) or state_cur(176) or state_cur(426) or state_cur(194) or state_cur(124) or state_cur(348) or ( state_cur(433) and in70 ) or ( state_cur(59) and not ( in16 ) ) or state_cur(87) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 0) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 0) ) or state_cur(10) or state_cur(465) or state_cur(21) or state_cur(136) or state_cur(135) or state_cur(171) or state_cur(354) or state_cur(183) or state_cur(96) or state_cur(317) or state_cur(122) or ( state_cur(80) and to_stdl(funccall2 = 2) ) or ( state_cur(79) and to_stdl(funccall2 = 2) ) or ( state_cur(64) and in17 ) or ( state_cur(64) and not ( in17 ) ) or ( state_cur(54) and not ( in15 ) ) or state_cur(430) or state_cur(52) or ( state_cur(45) and in12 ) or ( state_cur(45) and not ( in12 ) ) or ( state_cur(40) and not ( in10 ) ) or state_cur(188) or state_cur(38) or ( state_cur(121) and in26 ) or ( state_cur(454) and in76 ) or ( state_cur(17) and in3 ) or ( state_cur(82) and in24 ) or ( state_cur(396) and to_stdl(funccall0 = 15) ) or ( state_cur(396) and to_stdl(funccall0 = 16) ) or state_cur(140) or ( state_cur(252) and not ( in49 ) ) or state_cur(202) or ( state_cur(6) and in1 ) or ( state_cur(2) and in0 ) or ( state_cur(422) and in65 );
	out784_bufn <= state_cur(115) or state_cur(185);
	out3_bufn <= ( state_cur(419) and in64 ) or ( state_cur(278) and to_stdl(funccall9 = 0) ) or ( state_cur(278) and to_stdl(funccall9 = 1) ) or ( state_cur(439) and not ( in71 ) and to_stdl(funccall8 = 1) ) or ( state_cur(422) and in65 );
	out746_bufn <= state_cur(247) or state_cur(239) or state_cur(213) or state_cur(205);
	out528_bufn <= state_cur(297) or state_cur(332);
	out372_bufn <= state_cur(381) or state_cur(89);
	out418_bufn <= state_cur(334) or state_cur(299);
	out708_bufn <= state_cur(285) or state_cur(86);
	out706_bufn <= state_cur(193) or state_cur(362);
	out445_bufn <= state_cur(267) or state_cur(303);
	out1021_bufn <= state_cur(323) or state_cur(100);
	out405_bufn <= state_cur(193) or state_cur(115) or state_cur(312) or state_cur(311) or state_cur(310) or state_cur(95) or state_cur(185) or state_cur(176) or state_cur(362) or state_cur(194) or state_cur(348) or state_cur(96) or state_cur(317);
	out764_bufn <= state_cur(284) or state_cur(178);
	out581_bufn <= state_cur(253) or state_cur(133);
	out776_bufn <= state_cur(91) or state_cur(346);
	out213_bufn <= state_cur(184) or state_cur(154) or state_cur(255) or state_cur(12) or state_cur(68) or state_cur(63) or state_cur(57) or state_cur(50) or state_cur(49) or state_cur(44) or state_cur(42) or state_cur(34);
	out674_bufn <= state_cur(90) or state_cur(384);
	out1326_bufn <= state_cur(447) or state_cur(363) or ( state_cur(449) and in73 );
	out334_bufn <= ( state_cur(270) ) or ( state_cur(30) and in8 ) or ( state_cur(25) and in6 ) or ( state_cur(15) ) or ( state_cur(76) and in22 ) or ( state_cur(76) and not ( in22 ) ) or ( state_cur(74) and in21 );
	out843_bufn <= state_cur(275) or state_cur(165);
	out175_bufn <= state_cur(32) or state_cur(31) or ( state_cur(30) and not ( in8 ) );
	out1036_bufn <= state_cur(355) or state_cur(301);
	out1015_bufn <= state_cur(320) or state_cur(294);
	out236_bufn <= state_cur(378) or state_cur(429) or ( state_cur(427) and not ( in68 ) );
	out395_bufn <= ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 4) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 4) ) or state_cur(164) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 0) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 0) ) or state_cur(306);
	out1340_bufn <= state_cur(446) or state_cur(383) or ( state_cur(452) and in75 );
	out993_bufn <= state_cur(200) or state_cur(92);
	out356_bufn <= state_cur(149) or state_cur(302);
	out273_bufn <= state_cur(102) or state_cur(372);
	out403_bufn <= state_cur(176) or state_cur(317);
	out286_bufn <= state_cur(290) or state_cur(350);
	out364_bufn <= state_cur(176) or state_cur(194) or state_cur(124) or state_cur(348) or state_cur(87) or state_cur(354) or state_cur(183) or state_cur(122);
	out697_bufn <= state_cur(253) or state_cur(191) or ( state_cur(252) and in49 );
	out283_bufn <= state_cur(174) or state_cur(441) or ( state_cur(366) and not ( in53 ) );
	out282_bufn <= state_cur(331) or state_cur(56);
	out1319_bufn <= ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 3) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 3) ) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 2) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 2) ) or ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 1) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 1) );
	out409_bufn <= state_cur(326) or state_cur(296);
	out1092_bufn <= state_cur(339) or state_cur(155);
	out1075_bufn <= state_cur(356) or state_cur(95);
	out925_bufn <= ( state_cur(51) and to_stdl(funccall5 = 0) ) or ( state_cur(35) and to_stdl(funccall6 = 1) );
	out78_bufn <= state_cur(144) or state_cur(464) or state_cur(143) or state_cur(235) or state_cur(155) or state_cur(114) or state_cur(313) or state_cur(309) or state_cur(308) or state_cur(108) or state_cur(304) or state_cur(434) or state_cur(301) or state_cur(103) or state_cur(101) or state_cur(298) or state_cur(297) or state_cur(100) or state_cur(97) or state_cur(294) or state_cur(293) or state_cur(94) or state_cur(291) or state_cur(91) or state_cur(289) or state_cur(288) or state_cur(287) or state_cur(286) or state_cur(285) or state_cur(284) or state_cur(90) or state_cur(92) or state_cur(281) or state_cur(84) or state_cur(277) or state_cur(269) or state_cur(268) or state_cur(267) or state_cur(58) or state_cur(85) or state_cur(9) or state_cur(463) or state_cur(111) or state_cur(314) or state_cur(307) or state_cur(104) or state_cur(300) or state_cur(102) or state_cur(106) or state_cur(299) or state_cur(98) or state_cur(290) or state_cur(296) or state_cur(295) or state_cur(93) or state_cur(99) or state_cur(292) or state_cur(315) or state_cur(89) or state_cur(283) or state_cur(282) or state_cur(302) or state_cur(56) or state_cur(266) or state_cur(327);
	out1089_bufn <= state_cur(368) or state_cur(114);
	out362_bufn <= state_cur(124) or state_cur(87) or state_cur(171) or state_cur(354) or state_cur(183) or state_cur(122);
	out982_bufn <= state_cur(357) or state_cur(277);
	out979_bufn <= ( state_cur(82) and not ( in24 ) ) or state_cur(269);
	out952_bufn <= state_cur(113) or state_cur(268);
	out1109_bufn <= state_cur(464) or state_cur(177);
	out16_bufn <= state_cur(459) or state_cur(440) or state_cur(220) or state_cur(161) or state_cur(139) or state_cur(83) or state_cur(16) or state_cur(19) or state_cur(18) or state_cur(14) or state_cur(7) or state_cur(5) or state_cur(8) or state_cur(3);
	out703_bufn <= state_cur(310) or state_cur(362);
	out371_bufn <= state_cur(216) or state_cur(283);
	out956_bufn <= state_cur(271) or ( state_cur(256) ) or ( state_cur(254) );
	out1107_bufn <= state_cur(144) or state_cur(349);
	out1033_bufn <= state_cur(175) or state_cur(103);
	out148_bufn <= state_cur(146) or ( state_cur(121) and in26 );
	out351_bufn <= state_cur(321) or state_cur(223) or state_cur(224) or state_cur(107) or state_cur(83) or state_cur(16);
	out740_bufn <= ( state_cur(396) and to_stdl(funccall0 = 0) ) or ( state_cur(338) and in52 ) or ( state_cur(251) and in48 ) or ( state_cur(249) and not ( in47 ) ) or ( state_cur(249) and in47 ) or ( state_cur(246) and not ( in46 ) ) or ( state_cur(243) ) or ( state_cur(242) ) or ( state_cur(238) ) or ( state_cur(237) ) or ( state_cur(212) and in43 ) or ( state_cur(211) ) or ( state_cur(207) and to_stdl(funccall1 = 0) ) or ( state_cur(207) and to_stdl(funccall1 = 3) ) or ( state_cur(179) and in40 ) or ( state_cur(170) and in39 ) or ( state_cur(160) and in38 ) or ( state_cur(148) and in36 ) or ( state_cur(137) and not ( in34 ) ) or ( state_cur(130) and not ( in33 ) ) or ( state_cur(130) and in33 ) or ( state_cur(396) and to_stdl(funccall0 = 5) ) or ( state_cur(244) ) or ( state_cur(137) and in34 ) or ( state_cur(126) and not ( in32 ) and not ( in31 ) and not ( in30 ) and not ( in29 ) and in28 ) or ( state_cur(126) and not ( in32 ) and not ( in31 ) and not ( in30 ) and in29 ) or ( state_cur(126) and not ( in32 ) and not ( in31 ) and in30 ) or ( state_cur(126) and not ( in32 ) and in31 ) or state_cur(365);
	out391_bufn <= state_cur(127) or state_cur(4) or state_cur(425) or state_cur(306);
	out129_bufn <= state_cur(356) or ( state_cur(82) and in24 );
	out338_bufn <= ( state_cur(256) ) or ( state_cur(254) ) or ( state_cur(453) and to_stdl(funccall4 = 1) ) or ( state_cur(131) and to_stdl(funccall4 = 1) ) or ( state_cur(70) and to_stdl(funccall4 = 1) ) or state_cur(190) or state_cur(187) or state_cur(186) or ( state_cur(126) and in32 ) or ( state_cur(453) and to_stdl(funccall4 = 0) ) or ( state_cur(131) and to_stdl(funccall4 = 0) ) or ( state_cur(70) and to_stdl(funccall4 = 0) ) or state_cur(273) or ( state_cur(76) and in22 ) or ( state_cur(76) and not ( in22 ) );
	out425_bufn <= state_cur(55) or state_cur(300);
	out1078_bufn <= state_cur(311) or state_cur(310) or state_cur(95);
	out349_bufn <= ( state_cur(80) and to_stdl(funccall2 = 1) ) or ( state_cur(79) and to_stdl(funccall2 = 1) ) or ( state_cur(80) and to_stdl(funccall2 = 0) ) or ( state_cur(79) and to_stdl(funccall2 = 0) );
	out590_bufn <= state_cur(165) or state_cur(186) or ( state_cur(126) and in32 );
	out325_bufn <= state_cur(273) or state_cur(432) or state_cur(71) or ( state_cur(80) and to_stdl(funccall2 = 2) ) or ( state_cur(79) and to_stdl(funccall2 = 2) );
	out112_bufn <= state_cur(459) or state_cur(14) or state_cur(7) or state_cur(5);
	out224_bufn <= ( state_cur(54) and in15 ) or ( state_cur(53) and not ( in14 ) );
	out1220_bufn <= ( state_cur(265) and not ( not (in51) ) ) or ( state_cur(390) and not ( in54 ) );
	out1250_bufn <= ( state_cur(407) and in58 ) or ( state_cur(414) and in61 );
	out365_bufn <= ( state_cur(105) and in25 ) or state_cur(176) or state_cur(194) or state_cur(124) or state_cur(348) or state_cur(87) or state_cur(171) or state_cur(354) or state_cur(183) or state_cur(122);
	out699_bufn <= ( state_cur(453) and to_stdl(funccall4 = 1) ) or ( state_cur(131) and to_stdl(funccall4 = 1) ) or ( state_cur(70) and to_stdl(funccall4 = 1) ) or state_cur(191) or ( state_cur(252) and in49 );
	out488_bufn <= ( state_cur(105) and in25 ) or state_cur(171);
	out1069_bufn <= state_cur(404) or state_cur(108);
	out530_bufn <= state_cur(340) or state_cur(463);
	out326_bufn <= ( state_cur(452) and not ( in75 ) and to_stdl(funccall7 = 2) ) or ( state_cur(451) and not ( in74 ) and to_stdl(funccall7 = 2) ) or ( state_cur(80) and to_stdl(funccall2 = 2) ) or ( state_cur(79) and to_stdl(funccall2 = 2) );
	out602_bufn <= state_cur(255) or state_cur(12) or state_cur(163) or state_cur(11);
	out83_bufn <= state_cur(147) or state_cur(467) or state_cur(146) or state_cur(10) or state_cur(465) or state_cur(21) or state_cur(140);
	out311_bufn <= ( state_cur(433) and not ( in70 ) ) or ( state_cur(366) and in53 ) or state_cur(36) or state_cur(41) or ( state_cur(64) and in17 );
	out253_bufn <= state_cur(431) or ( state_cur(428) and not ( in69 ) ) or ( state_cur(427) and in68 ) or state_cur(426) or ( state_cur(45) and in12 );
	out209_bufn <= state_cur(426) or ( state_cur(39) and in9 );
	out1240_bufn <= ( state_cur(417) and in63 ) or state_cur(410) or ( state_cur(417) and not ( in63 ) ) or state_cur(398);
	out1018_bufn <= state_cur(325) or state_cur(97);
	out1152_bufn <= state_cur(429) or state_cur(441);
	out1236_bufn <= state_cur(408) or state_cur(406) or state_cur(405) or state_cur(402);
	out130_bufn <= state_cur(356) or state_cur(186) or ( state_cur(126) and in32 ) or ( state_cur(82) and in24 );
	out567_bufn <= ( state_cur(207) and to_stdl(funccall1 = 4) ) or ( state_cur(207) and to_stdl(funccall1 = 5) );
	out646_bufn <= ( state_cur(29) and in7 ) or ( state_cur(24) and in5 );

	-- Assignment of non-buffered outputs

	out26 <=
		state_cur(3);
	out2 <=
		state_cur(466) or state_cur(253) or state_cur(202) or state_cur(191) or state_cur(19) or state_cur(0);
	out931 <=
		state_cur(261);
	out715 <=
		state_cur(201);
	out410 <=
		state_cur(98);
	out628 <=
		state_cur(165);
	out734 <=
		state_cur(229) or state_cur(206);
	out942 <=
		state_cur(265);
	out122 <=
		state_cur(16);
	out892 <=
		state_cur(255);
	out601 <=
		state_cur(159);
	out809 <=
		state_cur(232);
	out376 <=
		state_cur(91);
	out241 <=
		state_cur(45);
	out986 <=
		state_cur(280);
	out1323 <=
		state_cur(446);
	out455 <=
		state_cur(117);
	out53 <=
		state_cur(377) or state_cur(354) or state_cur(306) or state_cur(305) or state_cur(140) or state_cur(4);
	out733 <=
		state_cur(206);
	out229 <=
		state_cur(41);
	out901 <=
		state_cur(469) or state_cur(462) or state_cur(461) or state_cur(445) or state_cur(257);
	out60 <=
		state_cur(425) or state_cur(377) or state_cur(306) or state_cur(305) or state_cur(127) or state_cur(4);
	out228 <=
		state_cur(444) or state_cur(441) or state_cur(430) or state_cur(68) or state_cur(67) or state_cur(57) or state_cur(41);
	out160 <=
		state_cur(25);
	out561 <=
		state_cur(150);
	out743 <=
		state_cur(208);
	out921 <=
		state_cur(259);
	out382 <=
		state_cur(93);
	out566 <=
		state_cur(151);
	out99 <=
		state_cur(255) or state_cur(163) or state_cur(12) or state_cur(11);
	out765 <=
		state_cur(217);
	out366 <=
		state_cur(88);
	out1005 <=
		state_cur(289);
	out1119 <=
		state_cur(345);
	out1356 <=
		state_cur(461);
	out25 <=
		state_cur(8) or state_cur(3);
	out802 <=
		state_cur(230);
	out918 <=
		state_cur(259) or state_cur(258);
	out258 <=
		state_cur(50);
	out640 <=
		state_cur(166);
	out710 <=
		state_cur(198);
	out1014 <=
		state_cur(294);
	out505 <=
		state_cur(443) or state_cur(437) or state_cur(133) or state_cur(132);
	out1303 <=
		state_cur(439);
	out424 <=
		state_cur(104);
	out920 <=
		state_cur(258);
	out180 <=
		state_cur(31);
	out974 <=
		state_cur(276);
	out1339 <=
		state_cur(450);
	out300 <=
		state_cur(64);
	out472 <=
		state_cur(123);
	out143 <=
		state_cur(324) or state_cur(20);
	out1301 <=
		state_cur(437);
	out479 <=
		state_cur(125);
	out464 <=
		state_cur(120);
	out643 <=
		state_cur(167);
	out636 <=
		state_cur(420) or state_cur(276) or state_cur(275) or state_cur(236) or state_cur(165);
	out1022 <=
		state_cur(297);
	out153 <=
		state_cur(23);
	out263 <=
		state_cur(51);
	out690 <=
		state_cur(213) or state_cur(187);
	out712 <=
		state_cur(199);
	out828 <=
		state_cur(235);
	out772 <=
		state_cur(220);
	out342 <=
		state_cur(76);
	out40 <=
		state_cur(465) or state_cur(425) or state_cur(306) or state_cur(127) or state_cur(87) or state_cur(4);
	out1223 <=
		state_cur(394);
	out443 <=
		state_cur(112);
	out679 <=
		state_cur(180);
	out1073 <=
		state_cur(309);
	out150 <=
		state_cur(21);
	out299 <=
		state_cur(68) or state_cur(63);
	out1349 <=
		state_cur(455);
	out1383 <=
		state_cur(471);
	out572 <=
		state_cur(153);
	out1298 <=
		state_cur(436);
	out1311 <=
		state_cur(442);
	out607 <=
		state_cur(161);
	out737 <=
		state_cur(207);
	out510 <=
		state_cur(396) or state_cur(365) or state_cur(207) or state_cur(134);
	out165 <=
		state_cur(28) or state_cur(26);
	out462 <=
		state_cur(119);
	out514 <=
		state_cur(136) or state_cur(135);
	out531 <=
		state_cur(143);
	out872 <=
		state_cur(243);
	out791 <=
		state_cur(226);
	out417 <=
		state_cur(101);
	out297 <=
		state_cur(63);
	out1121 <=
		state_cur(347);
	out614 <=
		state_cur(164);
	out64 <=
		state_cur(5);
	out589 <=
		state_cur(158);
	out231 <=
		state_cur(42);
	out888 <=
		state_cur(271) or state_cur(256) or state_cur(254);
	out1324 <=
		state_cur(447);
	out1150 <=
		state_cur(364);
	out1295 <=
		state_cur(435);
	out152 <=
		state_cur(159) or state_cur(22);
	out310 <=
		state_cur(444) or state_cur(67);
	out694 <=
		state_cur(189);
	out718 <=
		state_cur(202);
	out759 <=
		state_cur(214);
	out722 <=
		state_cur(203);
	out1387 <=
		state_cur(472);
	out82 <=
		state_cur(473) or state_cur(464) or state_cur(463) or state_cur(456) or state_cur(438) or state_cur(434) or state_cur(404) or state_cur(388) or
		state_cur(387) or state_cur(384) or state_cur(382) or state_cur(381) or state_cur(380) or state_cur(376) or state_cur(375) or state_cur(372) or
		state_cur(368) or state_cur(362) or state_cur(360) or state_cur(357) or state_cur(356) or state_cur(355) or state_cur(351) or state_cur(350) or
		state_cur(349) or state_cur(348) or state_cur(346) or state_cur(342) or state_cur(341) or state_cur(340) or state_cur(339) or state_cur(334) or
		state_cur(332) or state_cur(331) or state_cur(330) or state_cur(329) or state_cur(328) or state_cur(327) or state_cur(326) or state_cur(325) or
		state_cur(323) or state_cur(322) or state_cur(321) or state_cur(320) or state_cur(319) or state_cur(318) or state_cur(317) or state_cur(316) or
		state_cur(315) or state_cur(314) or state_cur(313) or state_cur(312) or state_cur(311) or state_cur(310) or state_cur(309) or state_cur(308) or
		state_cur(307) or state_cur(304) or state_cur(303) or state_cur(302) or state_cur(301) or state_cur(300) or state_cur(299) or state_cur(298) or
		state_cur(297) or state_cur(296) or state_cur(295) or state_cur(294) or state_cur(293) or state_cur(292) or state_cur(291) or state_cur(290) or
		state_cur(289) or state_cur(288) or state_cur(287) or state_cur(286) or state_cur(285) or state_cur(284) or state_cur(283) or state_cur(282) or
		state_cur(281) or state_cur(278) or state_cur(277) or state_cur(269) or state_cur(268) or state_cur(267) or state_cur(266) or state_cur(224) or
		state_cur(221) or state_cur(219) or state_cur(216) or state_cur(200) or state_cur(197) or state_cur(196) or state_cur(195) or state_cur(194) or
		state_cur(193) or state_cur(192) or state_cur(185) or state_cur(178) or state_cur(177) or state_cur(176) or state_cur(175) or state_cur(172) or
		state_cur(155) or state_cur(149) or state_cur(145) or state_cur(144) or state_cur(143) or state_cur(142) or state_cur(141) or state_cur(116) or
		state_cur(115) or state_cur(114) or state_cur(113) or state_cur(111) or state_cur(110) or state_cur(108) or state_cur(106) or state_cur(104) or
		state_cur(103) or state_cur(102) or state_cur(101) or state_cur(100) or state_cur(99) or state_cur(98) or state_cur(97) or state_cur(96) or
		state_cur(95) or state_cur(94) or state_cur(93) or state_cur(92) or state_cur(91) or state_cur(90) or state_cur(89) or state_cur(86) or
		state_cur(85) or state_cur(84) or state_cur(60) or state_cur(58) or state_cur(56) or state_cur(55) or state_cur(37) or state_cur(16) or
		state_cur(9);
	out1139 <=
		state_cur(361);
	out558 <=
		state_cur(147);
	out696 <=
		state_cur(190);
	out1381 <=
		state_cur(470);
	out1293 <=
		state_cur(435);
	out519 <=
		state_cur(139);
	out1292 <=
		state_cur(434);
	out895 <=
		state_cur(256);
	out1176 <=
		state_cur(429) or state_cur(379) or state_cur(378);
	out170 <=
		state_cur(173) or state_cur(27);
	out434 <=
		state_cur(109);
	out341 <=
		state_cur(77) or state_cur(75);
	out1007 <=
		state_cur(290);
	out595 <=
		state_cur(158);
	out874 <=
		state_cur(244);
	out1364 <=
		state_cur(464);
	out621 <=
		state_cur(164);
	out962 <=
		state_cur(273);
	out767 <=
		state_cur(374) or state_cur(220) or state_cur(217);
	out523 <=
		state_cur(139);
	out350 <=
		state_cur(81);
	out745 <=
		state_cur(209);
	out863 <=
		state_cur(241);
	out958 <=
		state_cur(272);
	out1182 <=
		state_cur(446) or state_cur(383);
	out13 <=
		state_cur(1);
	out1 <=
		state_cur(0);
	out1101 <=
		state_cur(336);
	out1344 <=
		state_cur(452);
	out749 <=
		state_cur(210);
	out972 <=
		state_cur(275);
	out289 <=
		state_cur(61);
	out1290 <=
		state_cur(432);
	out985 <=
		state_cur(279);
	out279 <=
		state_cur(57);
	out517 <=
		state_cur(138);
	out1035 <=
		state_cur(302);
	out1000 <=
		state_cur(287);
	out1085 <=
		state_cur(314);
	out1289 <=
		state_cur(431);
	out85 <=
		state_cur(377) or state_cur(305) or state_cur(124) or state_cur(10);
	out35 <=
		state_cur(306) or state_cur(183) or state_cur(171) or state_cur(147) or state_cur(146) or state_cur(4);
	out304 <=
		state_cur(65);
	out347 <=
		state_cur(80) or state_cur(79);
	out1190 <=
		state_cur(389);
	out649 <=
		state_cur(167);
	out156 <=
		state_cur(24);
	out1228 <=
		state_cur(396);
	out266 <=
		state_cur(51);
	out651 <=
		state_cur(168);
	out866 <=
		state_cur(242);
	out508 <=
		state_cur(133);
	out1114 <=
		state_cur(344);
	out245 <=
		state_cur(46);
	out44 <=
		state_cur(354) or state_cur(306) or state_cur(21) or state_cur(4);
	out1174 <=
		state_cur(431) or state_cur(378);
	out80 <=
		state_cur(9);
	out134 <=
		state_cur(17);
	out1187 <=
		state_cur(391) or state_cur(386);
	out1032 <=
		state_cur(301);
	out1287 <=
		state_cur(430);
	out989 <=
		state_cur(281);
	out538 <=
		state_cur(146);
	out1104 <=
		state_cur(337);
	out981 <=
		state_cur(278);
	out1286 <=
		state_cur(429);
	out724 <=
		state_cur(204);
	out487 <=
		state_cur(127);
	out658 <=
		state_cur(169);
	out1215 <=
		state_cur(393) or state_cur(390);
	out407 <=
		state_cur(97);
	out534 <=
		state_cur(144);
	out1175 <=
		state_cur(378);
	out858 <=
		state_cur(239);
	out1284 <=
		state_cur(429);
	out402 <=
		state_cur(356) or state_cur(171) or state_cur(146) or state_cur(95);
	out755 <=
		state_cur(212);
	out255 <=
		state_cur(48);
	out93 <=
		state_cur(11);
	out467 <=
		state_cur(122);
	out379 <=
		state_cur(92);
	out664 <=
		state_cur(174);
	out429 <=
		state_cur(106);
	out322 <=
		state_cur(123) or state_cur(81) or state_cur(71);
	out949 <=
		state_cur(268);
	out826 <=
		state_cur(389) or state_cur(235);
	out681 <=
		state_cur(181);
	out905 <=
		state_cur(462) or state_cur(461) or state_cur(445) or state_cur(257);
	out15 <=
		state_cur(2);
	out794 <=
		state_cur(227);
	out795 <=
		state_cur(228);
	out139 <=
		state_cur(19);
	out193 <=
		state_cur(35);
	out1019 <=
		state_cur(296);
	out171 <=
		state_cur(28);
	out173 <=
		state_cur(29);
	out610 <=
		state_cur(162);
	out1279 <=
		state_cur(427);
	out440 <=
		state_cur(111);
	out480 <=
		state_cur(134) or state_cur(125);
	out860 <=
		state_cur(239);
	out1158 <=
		state_cur(369);
	out189 <=
		state_cur(33);
	out902 <=
		state_cur(257);
	out1134 <=
		state_cur(358);
	out799 <=
		state_cur(229);
	out955 <=
		state_cur(270);
	out1278 <=
		state_cur(426);
	out1098 <=
		state_cur(335);
	out963 <=
		state_cur(274);
	out373 <=
		state_cur(90);
	out728 <=
		state_cur(213) or state_cur(205);
	out1160 <=
		state_cur(370);
	out570 <=
		state_cur(353) or state_cur(214) or state_cur(152);
	out937 <=
		state_cur(262);
	out1275 <=
		state_cur(426);
	out114 <=
		state_cur(14);
	out812 <=
		state_cur(233);
	out787 <=
		state_cur(225);
	out7 <=
		state_cur(421) or state_cur(420) or state_cur(415) or state_cur(413) or state_cur(412) or state_cur(408) or state_cur(406) or state_cur(405) or
		state_cur(402) or state_cur(401) or state_cur(275) or state_cur(261) or state_cur(165) or state_cur(0);
	out396 <=
		state_cur(95);
	out762 <=
		state_cur(215);
	out978 <=
		state_cur(277);
	out933 <=
		state_cur(410) or state_cur(398) or state_cur(261);
	out938 <=
		state_cur(263);
	out313 <=
		state_cur(67);
	out1131 <=
		state_cur(356);
	out778 <=
		state_cur(222);
	out848 <=
		state_cur(236);
	out882 <=
		state_cur(251) or state_cur(250) or state_cur(248);
	out1229 <=
		state_cur(398);
	out1180 <=
		state_cur(450) or state_cur(383);
	out1155 <=
		state_cur(367);
	out947 <=
		state_cur(267);
	out232 <=
		state_cur(426) or state_cur(258) or state_cur(158) or state_cur(42);
	out201 <=
		state_cur(36);
	out783 <=
		state_cur(223);
	out996 <=
		state_cur(284);
	out1094 <=
		state_cur(333);
	out420 <=
		state_cur(102);
	out107 <=
		state_cur(12);
	out1269 <=
		state_cur(425);
	out414 <=
		state_cur(100);
	out1011 <=
		state_cur(292);
	out333 <=
		state_cur(123) or state_cur(72);
	out296 <=
		state_cur(62);
	out335 <=
		state_cur(73);
	out726 <=
		state_cur(205);
	out1151 <=
		state_cur(366);
	out256 <=
		state_cur(49);
	out111 <=
		state_cur(255) or state_cur(12);
	out1068 <=
		state_cur(307);
	out202 <=
		state_cur(174) or state_cur(36);
	out1368 <=
		state_cur(467);
	out1181 <=
		state_cur(383);
	out1137 <=
		state_cur(359);
	out1308 <=
		state_cur(441);
	out768 <=
		state_cur(218);
	out500 <=
		state_cur(131);
	out14 <=
		state_cur(455) or state_cur(442) or state_cur(436) or state_cur(400) or state_cur(394) or state_cur(385) or state_cur(373) or state_cur(370) or
		state_cur(369) or state_cur(367) or state_cur(364) or state_cur(361) or state_cur(359) or state_cur(358) or state_cur(352) or state_cur(347) or
		state_cur(345) or state_cur(344) or state_cur(343) or state_cur(337) or state_cur(336) or state_cur(335) or state_cur(280) or state_cur(279) or
		state_cur(274) or state_cur(272) or state_cur(233) or state_cur(232) or state_cur(231) or state_cur(230) or state_cur(228) or state_cur(227) or
		state_cur(226) or state_cur(225) or state_cur(223) or state_cur(222) or state_cur(218) or state_cur(215) or state_cur(208) or state_cur(204) or
		state_cur(203) or state_cur(201) or state_cur(199) or state_cur(198) or state_cur(189) or state_cur(182) or state_cur(181) or state_cur(180) or
		state_cur(166) or state_cur(162) or state_cur(156) or state_cur(153) or state_cur(151) or state_cur(150) or state_cur(120) or state_cur(119) or
		state_cur(118) or state_cur(117) or state_cur(112) or state_cur(109) or state_cur(88) or state_cur(62) or state_cur(33) or state_cur(3) or
		state_cur(1);
	out1164 <=
		state_cur(371);
	out1125 <=
		state_cur(352);
	out1016 <=
		state_cur(295);
	out688 <=
		state_cur(186);
	out1026 <=
		state_cur(299);
	out1329 <=
		state_cur(449);
	out191 <=
		state_cur(34);
	out855 <=
		state_cur(238);
	out597 <=
		state_cur(258) or state_cur(158);
	out184 <=
		state_cur(32) or state_cur(31);
	out162 <=
		state_cur(26);
	out422 <=
		state_cur(103);
	out197 <=
		state_cur(188) or state_cur(38) or state_cur(35);
	out104 <=
		state_cur(12);
	out1266 <=
		state_cur(423);
	out117 <=
		state_cur(15);
	out1024 <=
		state_cur(298);
	out221 <=
		state_cur(41);
	out1088 <=
		state_cur(315);
	out1128 <=
		state_cur(354);
	out923 <=
		state_cur(260) or state_cur(259);
	out1029 <=
		state_cur(300);
	out137 <=
		state_cur(19) or state_cur(18);
	out515 <=
		state_cur(136);
	out991 <=
		state_cur(282);
	out1375 <=
		state_cur(468);
	out957 <=
		state_cur(271);
	out264 <=
		state_cur(430) or state_cur(52) or state_cur(51);
	out1262 <=
		state_cur(421);
	out663 <=
		state_cur(173);
	out1111 <=
		state_cur(343);
	out119 <=
		state_cur(15);
	out998 <=
		state_cur(286);
	out731 <=
		state_cur(206);
	out1366 <=
		state_cur(466);
	out320 <=
		state_cur(453) or state_cur(131) or state_cur(70);
	out208 <=
		state_cur(38);
	out994 <=
		state_cur(283);
	out136 <=
		state_cur(18);
	out1145 <=
		state_cur(363);
	out1126 <=
		state_cur(353);
	out478 <=
		state_cur(124);
	out753 <=
		state_cur(211);
	out1141 <=
		state_cur(362);
	out951 <=
		state_cur(269);
	out370 <=
		state_cur(89);
	out259 <=
		state_cur(57) or state_cur(50);
	out332 <=
		state_cur(72);
	out1370 <=
		state_cur(472) or state_cur(468);
	out281 <=
		state_cur(58);
	out234 <=
		state_cur(429) or state_cur(426) or state_cur(379) or state_cur(188) or state_cur(49) or state_cur(48) or state_cur(42);
	out314 <=
		state_cur(68);
	out1185 <=
		state_cur(385);
	out1353 <=
		state_cur(459);
	out907 <=
		state_cur(257);
	out1258 <=
		state_cur(420);
	out698 <=
		state_cur(191);
	out212 <=
		state_cur(40);
	out468 <=
		state_cur(467) or state_cur(377) or state_cur(305) or state_cur(122);
	out876 <=
		state_cur(245);
	out498 <=
		state_cur(129);
	out251 <=
		state_cur(379) or state_cur(48);
	out1009 <=
		state_cur(291);
	out656 <=
		state_cur(168);
	out612 <=
		state_cur(163);
	out177 <=
		state_cur(30);
	out944 <=
		state_cur(266);
	out894 <=
		state_cur(255);
	out928 <=
		state_cur(261) or state_cur(260);
	out267 <=
		state_cur(52);
	out384 <=
		state_cur(94);
	out1171 <=
		state_cur(374);
	out815 <=
		state_cur(234);
	out230 <=
		state_cur(260) or state_cur(259) or state_cur(57) or state_cur(41);
	out739 <=
		state_cur(365) or state_cur(207);
	out88 <=
		state_cur(467) or state_cur(465) or state_cur(425) or state_cur(354) or state_cur(348) or state_cur(317) or state_cur(312) or state_cur(311) or
		state_cur(310) or state_cur(194) or state_cur(193) or state_cur(185) or state_cur(183) or state_cur(176) or state_cur(171) or state_cur(147) or
		state_cur(146) or state_cur(140) or state_cur(127) or state_cur(124) or state_cur(122) or state_cur(115) or state_cur(96) or state_cur(87) or
		state_cur(21) or state_cur(10);
	out997 <=
		state_cur(285);
	out1362 <=
		state_cur(462);
	out806 <=
		state_cur(231);
	out1037 <=
		state_cur(304);
	out1147 <=
		state_cur(447) or state_cur(363);
	out1253 <=
		state_cur(471) or state_cur(470) or state_cur(458) or state_cur(418);
	out1169 <=
		state_cur(373);
	out316 <=
		state_cur(70);
	out317 <=
		state_cur(131) or state_cur(123) or state_cur(81) or state_cur(77) or state_cur(75) or state_cur(71) or state_cur(70);
	out133 <=
		state_cur(371) or state_cur(362) or state_cur(107) or state_cur(95) or state_cur(83) or state_cur(16);
	out1252 <=
		state_cur(418);
	out1096 <=
		state_cur(333);
	out186 <=
		state_cur(32);
	out1346 <=
		state_cur(453);
	out1146 <=
		state_cur(363);
	out363 <=
		state_cur(87);
	out887 <=
		state_cur(254);
	out659 <=
		state_cur(190) or state_cur(169);
	out661 <=
		state_cur(171);
	out346 <=
		state_cur(79);
	out270 <=
		state_cur(54);
	out1363 <=
		state_cur(463);
	out886 <=
		state_cur(253);
	out1341 <=
		state_cur(451);
	out92 <=
		state_cur(11);
	out1213 <=
		state_cur(390);
	out324 <=
		state_cur(71);
	out578 <=
		state_cur(156);
	out344 <=
		state_cur(77);
	out929 <=
		state_cur(260);
	out355 <=
		state_cur(84);
	out953 <=
		state_cur(270);
	out146 <=
		state_cur(324) or state_cur(261) or state_cur(20);
	out1365 <=
		state_cur(465);
	out348 <=
		state_cur(80);
	out358 <=
		state_cur(85);
	out513 <=
		state_cur(135);
	out1217 <=
		state_cur(391);
	out305 <=
		state_cur(67) or state_cur(65);
	out903 <=
		state_cur(461) or state_cur(257);
	out239 <=
		state_cur(44);
	out497 <=
		state_cur(134) or state_cur(129) or state_cur(128);
	out1337 <=
		state_cur(450);
	out861 <=
		state_cur(247) or state_cur(239);
	out448 <=
		state_cur(114);
	out1070 <=
		state_cur(308);
	out527 <=
		state_cur(140);
	out247 <=
		state_cur(47);
	out1091 <=
		state_cur(327);
	out496 <=
		state_cur(128);
	out328 <=
		state_cur(432) or state_cur(273) or state_cur(71);
	out1186 <=
		state_cur(386);
	out1309 <=
		state_cur(441);
	out526 <=
		state_cur(161) or state_cur(139);
	out199 <=
		state_cur(35);
	out154 <=
		state_cur(435) or state_cur(253) or state_cur(133) or state_cur(23);
	out1243 <=
		state_cur(410);
	out55 <=
		state_cur(377) or state_cur(306) or state_cur(305) or state_cur(4);
	out1082 <=
		state_cur(313);
	out240 <=
		state_cur(49) or state_cur(44);
	out1320 <=
		state_cur(445);
	out458 <=
		state_cur(118);
	out879 <=
		state_cur(247);
	out936 <=
		state_cur(264) or state_cur(263) or state_cur(262);
	out84 <=
		state_cur(10);
	out1221 <=
		state_cur(423) or state_cur(397) or state_cur(395) or state_cur(392);
	out1003 <=
		state_cur(288);
	out192 <=
		state_cur(42) or state_cur(34);
	out692 <=
		state_cur(188);
	out852 <=
		state_cur(237);
	out275 <=
		state_cur(56);
	out775 <=
		state_cur(440) or state_cur(220);
	out412 <=
		state_cur(99);
	out306 <=
		state_cur(66);
	out1013 <=
		state_cur(293);
	out1235 <=
		state_cur(400);
	out577 <=
		state_cur(184) or state_cur(163) or state_cur(154);
	out1166 <=
		state_cur(371);
	out432 <=
		state_cur(108);
	out1327 <=
		state_cur(448);
	out1378 <=
		state_cur(469);
	out49 <=
		state_cur(306) or state_cur(171) or state_cur(146) or state_cur(4);
	out65 <=
		state_cur(459) or state_cur(14) or state_cur(7) or state_cur(5);
	out246 <=
		state_cur(48) or state_cur(46);
	out939 <=
		state_cur(264);
	out504 <=
		state_cur(132);
	out667 <=
		state_cur(444) or state_cur(441) or state_cur(174);
	out683 <=
		state_cur(182);
	out686 <=
		state_cur(183);

	-- Assignment of buffered outputs

	out1057 <= out1057_buf;
	out59 <= out59_buf;
	out447 <= out447_buf;
	out157 <= out157_buf;
	out450 <= out450_buf;
	out1012 <= out1012_buf;
	out1072 <= out1072_buf;
	out999 <= out999_buf;
	out437 <= out437_buf;
	out415 <= out415_buf;
	out426 <= out426_buf;
	out375 <= out375_buf;
	out704 <= out704_buf;
	out973 <= out973_buf;
	out11 <= out11_buf;
	out549 <= out549_buf;
	out453 <= out453_buf;
	out1231 <= out1231_buf;
	out87 <= out87_buf;
	out401 <= out401_buf;
	out990 <= out990_buf;
	out378 <= out378_buf;
	out1302 <= out1302_buf;
	out27 <= out27_buf;
	out569 <= out569_buf;
	out1030 <= out1030_buf;
	out537 <= out537_buf;
	out77 <= out77_buf;
	out1318 <= out1318_buf;
	out533 <= out533_buf;
	out32 <= out32_buf;
	out1027 <= out1027_buf;
	out599 <= out599_buf;
	out668 <= out668_buf;
	out568 <= out568_buf;
	out225 <= out225_buf;
	out700 <= out700_buf;
	out638 <= out638_buf;
	out670 <= out670_buf;
	out433 <= out433_buf;
	out896 <= out896_buf;
	out575 <= out575_buf;
	out428 <= out428_buf;
	out72 <= out72_buf;
	out404 <= out404_buf;
	out98 <= out98_buf;
	out67 <= out67_buf;
	out635 <= out635_buf;
	out381 <= out381_buf;
	out222 <= out222_buf;
	out339 <= out339_buf;
	out268 <= out268_buf;
	out419 <= out419_buf;
	out559 <= out559_buf;
	out1002 <= out1002_buf;
	out1006 <= out1006_buf;
	out276 <= out276_buf;
	out205 <= out205_buf;
	out943 <= out943_buf;
	out1080 <= out1080_buf;
	out408 <= out408_buf;
	out252 <= out252_buf;
	out71 <= out71_buf;
	out672 <= out672_buf;
	out357 <= out357_buf;
	out441 <= out441_buf;
	out1084 <= out1084_buf;
	out144 <= out144_buf;
	out574 <= out574_buf;
	out210 <= out210_buf;
	out128 <= out128_buf;
	out360 <= out360_buf;
	out948 <= out948_buf;
	out506 <= out506_buf;
	out207 <= out207_buf;
	out1083 <= out1083_buf;
	out491 <= out491_buf;
	out4 <= out4_buf;
	out784 <= out784_buf;
	out3 <= out3_buf;
	out746 <= out746_buf;
	out528 <= out528_buf;
	out372 <= out372_buf;
	out418 <= out418_buf;
	out708 <= out708_buf;
	out706 <= out706_buf;
	out445 <= out445_buf;
	out1021 <= out1021_buf;
	out405 <= out405_buf;
	out764 <= out764_buf;
	out581 <= out581_buf;
	out776 <= out776_buf;
	out213 <= out213_buf;
	out674 <= out674_buf;
	out1326 <= out1326_buf;
	out334 <= out334_buf;
	out843 <= out843_buf;
	out175 <= out175_buf;
	out1036 <= out1036_buf;
	out1015 <= out1015_buf;
	out236 <= out236_buf;
	out395 <= out395_buf;
	out1340 <= out1340_buf;
	out993 <= out993_buf;
	out356 <= out356_buf;
	out273 <= out273_buf;
	out403 <= out403_buf;
	out286 <= out286_buf;
	out364 <= out364_buf;
	out697 <= out697_buf;
	out283 <= out283_buf;
	out282 <= out282_buf;
	out1319 <= out1319_buf;
	out409 <= out409_buf;
	out1092 <= out1092_buf;
	out1075 <= out1075_buf;
	out925 <= out925_buf;
	out78 <= out78_buf;
	out1089 <= out1089_buf;
	out362 <= out362_buf;
	out982 <= out982_buf;
	out979 <= out979_buf;
	out952 <= out952_buf;
	out1109 <= out1109_buf;
	out16 <= out16_buf;
	out703 <= out703_buf;
	out371 <= out371_buf;
	out956 <= out956_buf;
	out1107 <= out1107_buf;
	out1033 <= out1033_buf;
	out148 <= out148_buf;
	out351 <= out351_buf;
	out740 <= out740_buf;
	out391 <= out391_buf;
	out129 <= out129_buf;
	out338 <= out338_buf;
	out425 <= out425_buf;
	out1078 <= out1078_buf;
	out349 <= out349_buf;
	out590 <= out590_buf;
	out325 <= out325_buf;
	out112 <= out112_buf;
	out224 <= out224_buf;
	out1220 <= out1220_buf;
	out1250 <= out1250_buf;
	out365 <= out365_buf;
	out699 <= out699_buf;
	out488 <= out488_buf;
	out1069 <= out1069_buf;
	out530 <= out530_buf;
	out326 <= out326_buf;
	out602 <= out602_buf;
	out83 <= out83_buf;
	out311 <= out311_buf;
	out253 <= out253_buf;
	out209 <= out209_buf;
	out1240 <= out1240_buf;
	out1018 <= out1018_buf;
	out1152 <= out1152_buf;
	out1236 <= out1236_buf;
	out130 <= out130_buf;
	out567 <= out567_buf;
	out646 <= out646_buf;

end architecture;

