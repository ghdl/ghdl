package p is
  --  Comment
  type state_t is (s1, s2, s3);
end p;
