package pkg is
  component comp is
  end component;
end pkg;

entity comp is
end comp;
