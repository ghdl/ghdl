
-- Copyright (C) 1996 Morgan Kaufmann Publishers, Inc

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: ch_13_fg_13_24.vhd,v 1.1.1.1 2001-08-22 18:20:48 paw Exp $
-- $Revision: 1.1.1.1 $
--
-- ---------------------------------------------------------------------

configuration interlock_control_with_estimates of interlock_control is

  for detailed_timing

  end for;

  -- . . .

end configuration interlock_control_with_estimates;

--------------------------------------------------

configuration interlock_control_with_actual of interlock_control is

  for detailed_timing

    for ex_interlock_gate : nor_gate
      generic map ( Tpd01 => 320 ps, Tpd10 => 230 ps );
    end for;

    -- . . .

  end for;

end configuration interlock_control_with_actual;
