library ieee;use ieee.numeric_std.all;use ieee.std_logic_1164.all;entity t is
port(u:std'c;t:e(0);t:r(0));end;architecture t of t is type t is record
x:r range 0 to 0;end record;signal m:t;begin
t(((0)));f generic map(0);end architecture;