package function--
begin
X';