package function return of