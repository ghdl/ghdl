
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1750.vhd,v 1.2 2001-10-26 16:30:12 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c09s05b00x00p21n01i01750ent IS
  generic (g1: integer := 12);
  port (
    input1: in  bit ;
    input2: in  bit ;
    clk   : in  boolean;
    output: out bit);
END c09s05b00x00p21n01i01750ent;

ARCHITECTURE c09s05b00x00p21n01i01750arch OF c09s05b00x00p21n01i01750ent IS
  type boolvec is array (positive range <>) of boolean;
  function F (BB: boolvec) return boolean is
  begin
    return TRUE;
  end;
  
  signal i :  F boolean bus;
  signal k :  boolean ;
BEGIN
  i <= transport k;  -- Failure_here
  -- i is a guarded target while the statement is not a guarded assignment
  TESTING: PROCESS
  BEGIN
    assert FALSE 
      report "***FAILED TEST: c09s05b00x00p21n01i01750 - Ungarded signal can not assign to a guarded signal." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c09s05b00x00p21n01i01750arch;
