package mypkg is
  constant msg : string := "Message from mylib.mypkg";
end mypkg;
