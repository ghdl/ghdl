entity err is
end;

architecture behav of err is
  signal t2 : bit;
begin
  t0 <= '1';
end behav;
