package body gen1 is
  function get return natural is
  begin
    return v;
  end get;
end gen1;
