package pkga is
  constant a : natural := 5;
end;
