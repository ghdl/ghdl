entity t is end t;

architecture behav of t is
begin
  process
  begin
   report "val = " & "";
   wait;
  end process;
end;
