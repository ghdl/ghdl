package p is
  type state_t is
    (
      --  Comment
      s1,
      s2,
      s3);
end p;
