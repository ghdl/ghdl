architecture a2 of e2 is
  -- comments in design units (python doc-string style) :fail:
begin

end architecture;
