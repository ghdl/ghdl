LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE pkg IS
    TYPE test_record IS RECORD
        test : STD_LOGIC;
    END RECORD test_record;
END PACKAGE pkg;
