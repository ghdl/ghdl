entity ent is
end;

architecture a of ent is
    procedure p is
        type t is (A);
    begin
        for i in t loop
        end loop;
    end;
begin
end;
