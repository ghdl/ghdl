package package