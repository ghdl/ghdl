package float0generic0pkg is generic(package g is new I generic map(<>));--
function a(l:t;--
e:N:=0)--
return t;function m(r:e)return t;--
function t(g:d;--
h:h)return t;function p(s:t)return t;alias m is m;function r(e:t)return t;alias f is m;end float0generic0pkg;