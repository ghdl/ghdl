architecture arch of ent is
  signal b1 : bit;

  --  Comment for :b2:
  signal b2 : bit;
begin
end arch;
