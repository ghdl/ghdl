-- As packages define public elements like constants, types and sub-programs, we are intrested in such documentation too.:p2:
package p2 is
  -- comments in design units (python doc-string style):p2:
    -- might be multi line :p2:
end package;
