entity t is
end t1;
