library ieee;
use ieee.std_logic_1164.all;

entity top is
	port (
		clock : in  std_logic;
		reset : in  std_logic;
		start : in  std_logic;
		stdin_rdy : out std_logic;
		stdin_ack : in  std_logic;
		stdout_data : out std_logic_vector(31 downto 0);
		stdout_rdy : out std_logic;
		stdout_ack : in  std_logic;
		stdin_data : in  std_logic_vector(31 downto 0)
	);
end top;

architecture augh of top is

	-- Declaration of components

	component sub_147 is
		port (
			output : out std_logic_vector(63 downto 0);
			sign : in  std_logic;
			ge : out std_logic;
			in_a : in  std_logic_vector(63 downto 0);
			in_b : in  std_logic_vector(63 downto 0)
		);
	end component;

	component qq4_code4_table is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			ra0_addr : in  std_logic_vector(3 downto 0)
		);
	end component;

	component qq6_code6_table is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			ra0_addr : in  std_logic_vector(5 downto 0)
		);
	end component;

	component wl_code_table is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			ra0_addr : in  std_logic_vector(3 downto 0)
		);
	end component;

	component ilb_table is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			ra0_addr : in  std_logic_vector(4 downto 0)
		);
	end component;

	component decis_levl is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			ra0_addr : in  std_logic_vector(4 downto 0)
		);
	end component;

	component quant26bt_pos is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			ra0_addr : in  std_logic_vector(4 downto 0)
		);
	end component;

	component quant26bt_neg is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			ra0_addr : in  std_logic_vector(4 downto 0)
		);
	end component;

	component qq2_code2_table is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			ra0_addr : in  std_logic_vector(1 downto 0)
		);
	end component;

	component wh_code_table is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			ra0_addr : in  std_logic_vector(1 downto 0)
		);
	end component;

	component cmp_694 is
		port (
			in1 : in  std_logic_vector(31 downto 0);
			in0 : in  std_logic_vector(31 downto 0);
			eq : out std_logic
		);
	end component;

	component cmp_700 is
		port (
			in1 : in  std_logic_vector(31 downto 0);
			in0 : in  std_logic_vector(31 downto 0);
			eq : out std_logic
		);
	end component;

	component sub_144 is
		port (
			output : out std_logic_vector(63 downto 0);
			le : out std_logic;
			sign : in  std_logic;
			ge : out std_logic;
			in_a : in  std_logic_vector(63 downto 0);
			in_b : in  std_logic_vector(63 downto 0)
		);
	end component;

	component mul_145 is
		port (
			output : out std_logic_vector(63 downto 0);
			in_a : in  std_logic_vector(63 downto 0);
			in_b : in  std_logic_vector(31 downto 0)
		);
	end component;

	component mul_146 is
		port (
			output : out std_logic_vector(63 downto 0);
			in_a : in  std_logic_vector(63 downto 0);
			in_b : in  std_logic_vector(31 downto 0)
		);
	end component;

	component sub_143 is
		port (
			output : out std_logic_vector(63 downto 0);
			lt : out std_logic;
			le : out std_logic;
			sign : in  std_logic;
			gt : out std_logic;
			in_a : in  std_logic_vector(63 downto 0);
			in_b : in  std_logic_vector(63 downto 0)
		);
	end component;

	component add_142 is
		port (
			output : out std_logic_vector(63 downto 0);
			in_a : in  std_logic_vector(63 downto 0);
			in_b : in  std_logic_vector(63 downto 0)
		);
	end component;

	component test_data is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			wa0_addr : in  std_logic_vector(6 downto 0);
			wa0_en : in  std_logic;
			ra0_addr : in  std_logic_vector(6 downto 0);
			wa0_data : in  std_logic_vector(31 downto 0);
			ra1_data : out std_logic_vector(31 downto 0);
			ra1_addr : in  std_logic_vector(6 downto 0)
		);
	end component;

	component shr_141 is
		port (
			output : out std_logic_vector(31 downto 0);
			input : in  std_logic_vector(31 downto 0);
			shift : in  std_logic_vector(5 downto 0);
			padding : in  std_logic
		);
	end component;

	component compressed is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			wa0_addr : in  std_logic_vector(6 downto 0);
			wa0_en : in  std_logic;
			ra0_addr : in  std_logic_vector(6 downto 0);
			wa0_data : in  std_logic_vector(31 downto 0)
		);
	end component;

	component result is
		port (
			clk : in  std_logic;
			ra0_data : out std_logic_vector(31 downto 0);
			wa0_addr : in  std_logic_vector(6 downto 0);
			wa0_en : in  std_logic;
			ra0_addr : in  std_logic_vector(6 downto 0);
			wa0_data : in  std_logic_vector(31 downto 0)
		);
	end component;

	component cmp_662 is
		port (
			in1 : in  std_logic_vector(31 downto 0);
			in0 : in  std_logic_vector(31 downto 0);
			eq : out std_logic
		);
	end component;

	component cmp_673 is
		port (
			in1 : in  std_logic_vector(31 downto 0);
			in0 : in  std_logic_vector(31 downto 0);
			eq : out std_logic
		);
	end component;

	component mul_148 is
		port (
			output : out std_logic_vector(63 downto 0);
			in_a : in  std_logic_vector(32 downto 0);
			in_b : in  std_logic_vector(31 downto 0)
		);
	end component;

	component mul_149 is
		port (
			output : out std_logic_vector(63 downto 0);
			in_a : in  std_logic_vector(32 downto 0);
			in_b : in  std_logic_vector(31 downto 0)
		);
	end component;

	component add_153 is
		port (
			output : out std_logic_vector(63 downto 0);
			in_a : in  std_logic_vector(63 downto 0);
			in_b : in  std_logic_vector(63 downto 0)
		);
	end component;

	component add_154 is
		port (
			output : out std_logic_vector(63 downto 0);
			in_a : in  std_logic_vector(63 downto 0);
			in_b : in  std_logic_vector(63 downto 0)
		);
	end component;

	component add_155 is
		port (
			output : out std_logic_vector(63 downto 0);
			in_a : in  std_logic_vector(63 downto 0);
			in_b : in  std_logic_vector(63 downto 0)
		);
	end component;

	component mul_156 is
		port (
			output : out std_logic_vector(63 downto 0);
			in_a : in  std_logic_vector(32 downto 0);
			in_b : in  std_logic_vector(31 downto 0)
		);
	end component;

	component add_159 is
		port (
			output : out std_logic_vector(31 downto 0);
			in_a : in  std_logic_vector(31 downto 0);
			in_b : in  std_logic_vector(31 downto 0)
		);
	end component;

	component sub_160 is
		port (
			output : out std_logic_vector(63 downto 0);
			lt : out std_logic;
			le : out std_logic;
			sign : in  std_logic;
			ge : out std_logic;
			in_a : in  std_logic_vector(63 downto 0);
			in_b : in  std_logic_vector(63 downto 0)
		);
	end component;

	component mul_161 is
		port (
			output : out std_logic_vector(63 downto 0);
			in_a : in  std_logic_vector(32 downto 0);
			in_b : in  std_logic_vector(31 downto 0)
		);
	end component;

	component fsm_163 is
		port (
			clock : in  std_logic;
			reset : in  std_logic;
			out91 : out std_logic;
			out92 : out std_logic;
			out93 : out std_logic;
			in7 : in  std_logic;
			out94 : out std_logic;
			out95 : out std_logic;
			out98 : out std_logic;
			out100 : out std_logic;
			out101 : out std_logic;
			out102 : out std_logic;
			out104 : out std_logic;
			out105 : out std_logic;
			out106 : out std_logic;
			out107 : out std_logic;
			out108 : out std_logic;
			out109 : out std_logic;
			out111 : out std_logic;
			out114 : out std_logic;
			out116 : out std_logic;
			out118 : out std_logic;
			out119 : out std_logic;
			out120 : out std_logic;
			out128 : out std_logic;
			out130 : out std_logic;
			out131 : out std_logic;
			out132 : out std_logic;
			out137 : out std_logic;
			in8 : in  std_logic;
			out152 : out std_logic;
			out155 : out std_logic;
			out156 : out std_logic;
			out31 : out std_logic;
			in2 : in  std_logic;
			out28 : out std_logic;
			out29 : out std_logic;
			out30 : out std_logic;
			out26 : out std_logic;
			out27 : out std_logic;
			out24 : out std_logic;
			out25 : out std_logic;
			out77 : out std_logic;
			out79 : out std_logic;
			out80 : out std_logic;
			out82 : out std_logic;
			out34 : out std_logic;
			out35 : out std_logic;
			out36 : out std_logic;
			out32 : out std_logic;
			out33 : out std_logic;
			out40 : out std_logic;
			out41 : out std_logic;
			out88 : out std_logic;
			out89 : out std_logic;
			out21 : out std_logic;
			out22 : out std_logic;
			out23 : out std_logic;
			out73 : out std_logic;
			out76 : out std_logic;
			in6 : in  std_logic;
			out70 : out std_logic;
			out12 : out std_logic;
			out13 : out std_logic;
			out14 : out std_logic;
			out17 : out std_logic;
			out18 : out std_logic;
			out19 : out std_logic;
			out20 : out std_logic;
			out9 : out std_logic;
			out11 : out std_logic;
			out8 : out std_logic;
			out2 : out std_logic;
			out4 : out std_logic;
			out5 : out std_logic;
			in1 : in  std_logic;
			out6 : out std_logic;
			out7 : out std_logic;
			out0 : out std_logic;
			out1 : out std_logic;
			out37 : out std_logic;
			out38 : out std_logic;
			out39 : out std_logic;
			out1222 : out std_logic;
			out1223 : out std_logic;
			out1224 : out std_logic;
			out1225 : out std_logic;
			out1226 : out std_logic;
			out1228 : out std_logic;
			out1230 : out std_logic;
			in0 : in  std_logic;
			out67 : out std_logic;
			out68 : out std_logic;
			out65 : out std_logic;
			out66 : out std_logic;
			in5 : in  std_logic;
			out62 : out std_logic;
			out58 : out std_logic;
			out56 : out std_logic;
			in4 : in  std_logic;
			out57 : out std_logic;
			out54 : out std_logic;
			out55 : out std_logic;
			out51 : out std_logic;
			out52 : out std_logic;
			out53 : out std_logic;
			in3 : in  std_logic;
			out46 : out std_logic;
			out47 : out std_logic;
			out48 : out std_logic;
			out49 : out std_logic;
			out50 : out std_logic;
			out42 : out std_logic;
			out43 : out std_logic;
			out44 : out std_logic;
			out45 : out std_logic;
			in9 : in  std_logic;
			in10 : in  std_logic;
			out171 : out std_logic;
			in11 : in  std_logic;
			out191 : out std_logic;
			out207 : out std_logic;
			out208 : out std_logic;
			out209 : out std_logic;
			out212 : out std_logic;
			out213 : out std_logic;
			out216 : out std_logic;
			out220 : out std_logic;
			out221 : out std_logic;
			out223 : out std_logic;
			out224 : out std_logic;
			out226 : out std_logic;
			out227 : out std_logic;
			out228 : out std_logic;
			out229 : out std_logic;
			out230 : out std_logic;
			out233 : out std_logic;
			out235 : out std_logic;
			out236 : out std_logic;
			out237 : out std_logic;
			out238 : out std_logic;
			out239 : out std_logic;
			out241 : out std_logic;
			out250 : out std_logic;
			out258 : out std_logic;
			out259 : out std_logic;
			out261 : out std_logic;
			out270 : out std_logic;
			out276 : out std_logic;
			out277 : out std_logic;
			out283 : out std_logic;
			out285 : out std_logic;
			out287 : out std_logic;
			out290 : out std_logic;
			out291 : out std_logic;
			out293 : out std_logic;
			out301 : out std_logic;
			out303 : out std_logic;
			out304 : out std_logic;
			out315 : out std_logic;
			out319 : out std_logic;
			out321 : out std_logic;
			out330 : out std_logic;
			out335 : out std_logic;
			out338 : out std_logic;
			out341 : out std_logic;
			out342 : out std_logic;
			out344 : out std_logic;
			out347 : out std_logic;
			out351 : out std_logic;
			out354 : out std_logic;
			out355 : out std_logic;
			out356 : out std_logic;
			out357 : out std_logic;
			out358 : out std_logic;
			out360 : out std_logic;
			out361 : out std_logic;
			out362 : out std_logic;
			out365 : out std_logic;
			out367 : out std_logic;
			out368 : out std_logic;
			out370 : out std_logic;
			out375 : out std_logic;
			out376 : out std_logic;
			out378 : out std_logic;
			out381 : out std_logic;
			out382 : out std_logic;
			out386 : out std_logic;
			out387 : out std_logic;
			out388 : out std_logic;
			out390 : out std_logic;
			out392 : out std_logic;
			out393 : out std_logic;
			out394 : out std_logic;
			out397 : out std_logic;
			out403 : out std_logic;
			out404 : out std_logic;
			out408 : out std_logic;
			out409 : out std_logic;
			out410 : out std_logic;
			out412 : out std_logic;
			out416 : out std_logic;
			out417 : out std_logic;
			out418 : out std_logic;
			out419 : out std_logic;
			out420 : out std_logic;
			out421 : out std_logic;
			out424 : out std_logic;
			out425 : out std_logic;
			out430 : out std_logic;
			out431 : out std_logic;
			out434 : out std_logic;
			out436 : out std_logic;
			out438 : out std_logic;
			out439 : out std_logic;
			out440 : out std_logic;
			out441 : out std_logic;
			out442 : out std_logic;
			out443 : out std_logic;
			out444 : out std_logic;
			out445 : out std_logic;
			out446 : out std_logic;
			out447 : out std_logic;
			out448 : out std_logic;
			out450 : out std_logic;
			out451 : out std_logic;
			out454 : out std_logic;
			out457 : out std_logic;
			out460 : out std_logic;
			out463 : out std_logic;
			out465 : out std_logic;
			out466 : out std_logic;
			out472 : out std_logic;
			out473 : out std_logic;
			out475 : out std_logic;
			out476 : out std_logic;
			out479 : out std_logic;
			out480 : out std_logic;
			out481 : out std_logic;
			out482 : out std_logic;
			out484 : out std_logic;
			out485 : out std_logic;
			out489 : out std_logic;
			out491 : out std_logic;
			out494 : out std_logic;
			out497 : out std_logic;
			out500 : out std_logic;
			out503 : out std_logic;
			out504 : out std_logic;
			out505 : out std_logic;
			out508 : out std_logic;
			out509 : out std_logic;
			out513 : out std_logic;
			out514 : out std_logic;
			out516 : out std_logic;
			out521 : out std_logic;
			out523 : out std_logic;
			out524 : out std_logic;
			out525 : out std_logic;
			out530 : out std_logic;
			out532 : out std_logic;
			out533 : out std_logic;
			out535 : out std_logic;
			out536 : out std_logic;
			out539 : out std_logic;
			out541 : out std_logic;
			out543 : out std_logic;
			out545 : out std_logic;
			out547 : out std_logic;
			out549 : out std_logic;
			out550 : out std_logic;
			out552 : out std_logic;
			out558 : out std_logic;
			out559 : out std_logic;
			out563 : out std_logic;
			out566 : out std_logic;
			out572 : out std_logic;
			out573 : out std_logic;
			out576 : out std_logic;
			out577 : out std_logic;
			out581 : out std_logic;
			out582 : out std_logic;
			out590 : out std_logic;
			out591 : out std_logic;
			out592 : out std_logic;
			out593 : out std_logic;
			out595 : out std_logic;
			out611 : out std_logic;
			out619 : out std_logic;
			out638 : out std_logic;
			out643 : out std_logic;
			out644 : out std_logic;
			out645 : out std_logic;
			out646 : out std_logic;
			out648 : out std_logic;
			out650 : out std_logic;
			out652 : out std_logic;
			out657 : out std_logic;
			out659 : out std_logic;
			out662 : out std_logic;
			out677 : out std_logic;
			out678 : out std_logic;
			out679 : out std_logic;
			out680 : out std_logic;
			out682 : out std_logic;
			out686 : out std_logic;
			out692 : out std_logic;
			out1218 : out std_logic;
			out1219 : out std_logic;
			out1220 : out std_logic;
			out1221 : out std_logic;
			out695 : out std_logic;
			out697 : out std_logic;
			out706 : out std_logic;
			out719 : out std_logic;
			out729 : out std_logic;
			out744 : out std_logic;
			out746 : out std_logic;
			out748 : out std_logic;
			out833 : out std_logic;
			out834 : out std_logic;
			out836 : out std_logic;
			out837 : out std_logic;
			out839 : out std_logic;
			out840 : out std_logic;
			out841 : out std_logic;
			out844 : out std_logic;
			out845 : out std_logic;
			out846 : out std_logic;
			out848 : out std_logic;
			out850 : out std_logic;
			out852 : out std_logic;
			out854 : out std_logic;
			out856 : out std_logic;
			out858 : out std_logic;
			out860 : out std_logic;
			out863 : out std_logic;
			out865 : out std_logic;
			out866 : out std_logic;
			out873 : out std_logic;
			out877 : out std_logic;
			out888 : out std_logic;
			out891 : out std_logic;
			out893 : out std_logic;
			out895 : out std_logic;
			out898 : out std_logic;
			out900 : out std_logic;
			out902 : out std_logic;
			out903 : out std_logic;
			out904 : out std_logic;
			out905 : out std_logic;
			out906 : out std_logic;
			out907 : out std_logic;
			out908 : out std_logic;
			out909 : out std_logic;
			out910 : out std_logic;
			out912 : out std_logic;
			out913 : out std_logic;
			out914 : out std_logic;
			out915 : out std_logic;
			out917 : out std_logic;
			out920 : out std_logic;
			out921 : out std_logic;
			out924 : out std_logic;
			out934 : out std_logic;
			out935 : out std_logic;
			out937 : out std_logic;
			out938 : out std_logic;
			out940 : out std_logic;
			out943 : out std_logic;
			out945 : out std_logic;
			out957 : out std_logic;
			out958 : out std_logic;
			out962 : out std_logic;
			out968 : out std_logic;
			out972 : out std_logic;
			out973 : out std_logic;
			out974 : out std_logic;
			out975 : out std_logic;
			out976 : out std_logic;
			out980 : out std_logic;
			out986 : out std_logic;
			out988 : out std_logic;
			out989 : out std_logic;
			out990 : out std_logic;
			out1004 : out std_logic;
			out1008 : out std_logic;
			out999 : out std_logic;
			out1000 : out std_logic;
			out1002 : out std_logic;
			out1003 : out std_logic;
			out1050 : out std_logic;
			out1052 : out std_logic;
			out1053 : out std_logic;
			out1055 : out std_logic;
			out1056 : out std_logic;
			out1057 : out std_logic;
			out1059 : out std_logic;
			out1015 : out std_logic;
			out1025 : out std_logic;
			out1026 : out std_logic;
			out1038 : out std_logic;
			out1039 : out std_logic;
			out1042 : out std_logic;
			out1043 : out std_logic;
			out1046 : out std_logic;
			out1048 : out std_logic;
			out1061 : out std_logic;
			out1063 : out std_logic;
			out1064 : out std_logic;
			out1067 : out std_logic;
			out1068 : out std_logic;
			out1069 : out std_logic;
			out1071 : out std_logic;
			out1073 : out std_logic;
			out1076 : out std_logic;
			out1077 : out std_logic;
			out1078 : out std_logic;
			out1080 : out std_logic;
			out1081 : out std_logic;
			out1083 : out std_logic;
			out1085 : out std_logic;
			out1087 : out std_logic;
			out1089 : out std_logic;
			out1092 : out std_logic;
			out1096 : out std_logic;
			out1100 : out std_logic;
			out1103 : out std_logic;
			out1115 : out std_logic;
			out1122 : out std_logic;
			out1123 : out std_logic;
			out1127 : out std_logic;
			out1130 : out std_logic;
			out1133 : out std_logic;
			out1138 : out std_logic;
			out1139 : out std_logic;
			out1140 : out std_logic;
			out1141 : out std_logic;
			out1142 : out std_logic;
			out1143 : out std_logic;
			out1144 : out std_logic;
			out1145 : out std_logic;
			out1146 : out std_logic;
			out1147 : out std_logic;
			out1148 : out std_logic;
			out1149 : out std_logic;
			out1150 : out std_logic;
			out1151 : out std_logic;
			out1152 : out std_logic;
			out1153 : out std_logic;
			out1154 : out std_logic;
			out1155 : out std_logic;
			out1156 : out std_logic;
			out1157 : out std_logic;
			out1158 : out std_logic;
			out1159 : out std_logic;
			out1160 : out std_logic;
			out1161 : out std_logic;
			out1162 : out std_logic;
			out1163 : out std_logic;
			out1164 : out std_logic;
			out1165 : out std_logic;
			out1166 : out std_logic;
			out1167 : out std_logic;
			out1168 : out std_logic;
			out1169 : out std_logic;
			out1170 : out std_logic;
			out1171 : out std_logic;
			out1172 : out std_logic;
			out1173 : out std_logic;
			out1174 : out std_logic;
			out1175 : out std_logic;
			out1176 : out std_logic;
			out1177 : out std_logic;
			out1178 : out std_logic;
			out1179 : out std_logic;
			out1180 : out std_logic;
			out1181 : out std_logic;
			out1182 : out std_logic;
			out1183 : out std_logic;
			out1184 : out std_logic;
			out1185 : out std_logic;
			out1186 : out std_logic;
			out1187 : out std_logic;
			out1188 : out std_logic;
			out1189 : out std_logic;
			out1190 : out std_logic;
			out1191 : out std_logic;
			out1192 : out std_logic;
			out1193 : out std_logic;
			out1194 : out std_logic;
			out1195 : out std_logic;
			out1196 : out std_logic;
			out1197 : out std_logic;
			out1198 : out std_logic;
			out1199 : out std_logic;
			out1200 : out std_logic;
			out1201 : out std_logic;
			out1202 : out std_logic;
			out1203 : out std_logic;
			out1204 : out std_logic;
			out1205 : out std_logic;
			out1206 : out std_logic;
			out1207 : out std_logic;
			out1208 : out std_logic;
			out1209 : out std_logic;
			out1210 : out std_logic;
			out1211 : out std_logic;
			out1212 : out std_logic;
			out1213 : out std_logic;
			out1214 : out std_logic;
			out1215 : out std_logic;
			out1216 : out std_logic;
			out1217 : out std_logic
		);
	end component;

	-- Declaration of signals

	signal sig_clock : std_logic;
	signal sig_reset : std_logic;
	signal augh_test_23 : std_logic;
	signal augh_test_24 : std_logic;
	signal augh_test_78 : std_logic;
	signal augh_test_92 : std_logic;
	signal sig_start : std_logic;
	signal augh_test_113 : std_logic;
	signal augh_test_124 : std_logic;
	signal augh_test_135 : std_logic;
	signal augh_test_137 : std_logic;
	signal augh_test_138 : std_logic;
	signal sig_782 : std_logic;
	signal sig_783 : std_logic;
	signal sig_784 : std_logic;
	signal sig_785 : std_logic;
	signal sig_786 : std_logic;
	signal sig_787 : std_logic;
	signal sig_788 : std_logic;
	signal sig_789 : std_logic;
	signal sig_790 : std_logic;
	signal sig_791 : std_logic;
	signal sig_792 : std_logic;
	signal sig_793 : std_logic;
	signal sig_794 : std_logic;
	signal sig_795 : std_logic;
	signal sig_796 : std_logic;
	signal sig_797 : std_logic;
	signal sig_798 : std_logic;
	signal sig_799 : std_logic;
	signal sig_800 : std_logic;
	signal sig_801 : std_logic;
	signal sig_802 : std_logic;
	signal sig_803 : std_logic;
	signal sig_804 : std_logic;
	signal sig_805 : std_logic;
	signal sig_806 : std_logic;
	signal sig_807 : std_logic;
	signal sig_808 : std_logic;
	signal sig_809 : std_logic;
	signal sig_810 : std_logic;
	signal sig_811 : std_logic;
	signal sig_812 : std_logic;
	signal sig_813 : std_logic;
	signal sig_814 : std_logic;
	signal sig_815 : std_logic;
	signal sig_816 : std_logic;
	signal sig_817 : std_logic;
	signal sig_818 : std_logic;
	signal sig_819 : std_logic;
	signal sig_820 : std_logic;
	signal sig_821 : std_logic;
	signal sig_822 : std_logic;
	signal sig_823 : std_logic;
	signal sig_824 : std_logic;
	signal sig_825 : std_logic;
	signal sig_826 : std_logic;
	signal sig_827 : std_logic;
	signal sig_828 : std_logic;
	signal sig_829 : std_logic;
	signal sig_830 : std_logic;
	signal sig_831 : std_logic;
	signal sig_832 : std_logic;
	signal sig_833 : std_logic;
	signal sig_834 : std_logic;
	signal sig_835 : std_logic;
	signal sig_836 : std_logic;
	signal sig_837 : std_logic;
	signal sig_838 : std_logic;
	signal sig_839 : std_logic;
	signal sig_840 : std_logic;
	signal sig_841 : std_logic;
	signal sig_842 : std_logic;
	signal sig_843 : std_logic;
	signal sig_844 : std_logic;
	signal sig_845 : std_logic;
	signal sig_846 : std_logic;
	signal sig_847 : std_logic;
	signal sig_848 : std_logic;
	signal sig_849 : std_logic;
	signal sig_850 : std_logic;
	signal sig_851 : std_logic;
	signal sig_852 : std_logic;
	signal sig_853 : std_logic;
	signal sig_854 : std_logic;
	signal sig_855 : std_logic;
	signal sig_856 : std_logic;
	signal sig_857 : std_logic;
	signal sig_858 : std_logic;
	signal sig_859 : std_logic;
	signal sig_860 : std_logic;
	signal sig_861 : std_logic;
	signal sig_862 : std_logic;
	signal sig_863 : std_logic;
	signal sig_864 : std_logic;
	signal sig_865 : std_logic;
	signal sig_866 : std_logic;
	signal sig_867 : std_logic;
	signal sig_868 : std_logic;
	signal sig_869 : std_logic;
	signal sig_870 : std_logic;
	signal sig_871 : std_logic;
	signal sig_872 : std_logic;
	signal sig_873 : std_logic;
	signal sig_874 : std_logic;
	signal sig_875 : std_logic;
	signal sig_876 : std_logic;
	signal sig_877 : std_logic;
	signal sig_878 : std_logic;
	signal sig_879 : std_logic;
	signal sig_880 : std_logic;
	signal sig_881 : std_logic;
	signal sig_882 : std_logic;
	signal sig_883 : std_logic;
	signal sig_884 : std_logic;
	signal sig_885 : std_logic;
	signal sig_886 : std_logic;
	signal sig_887 : std_logic;
	signal sig_888 : std_logic;
	signal sig_889 : std_logic;
	signal sig_890 : std_logic;
	signal sig_891 : std_logic;
	signal sig_892 : std_logic;
	signal sig_893 : std_logic;
	signal sig_894 : std_logic;
	signal sig_895 : std_logic;
	signal sig_896 : std_logic;
	signal sig_897 : std_logic;
	signal sig_898 : std_logic;
	signal sig_899 : std_logic;
	signal sig_900 : std_logic;
	signal sig_901 : std_logic;
	signal sig_902 : std_logic;
	signal sig_903 : std_logic;
	signal sig_904 : std_logic;
	signal sig_905 : std_logic;
	signal sig_906 : std_logic;
	signal sig_907 : std_logic;
	signal sig_908 : std_logic;
	signal sig_909 : std_logic;
	signal sig_910 : std_logic;
	signal sig_911 : std_logic;
	signal sig_912 : std_logic;
	signal sig_913 : std_logic;
	signal sig_914 : std_logic;
	signal sig_915 : std_logic;
	signal sig_916 : std_logic;
	signal sig_917 : std_logic;
	signal sig_918 : std_logic;
	signal sig_919 : std_logic;
	signal sig_920 : std_logic;
	signal sig_921 : std_logic;
	signal sig_922 : std_logic;
	signal sig_923 : std_logic;
	signal sig_924 : std_logic;
	signal sig_925 : std_logic;
	signal sig_926 : std_logic;
	signal sig_927 : std_logic;
	signal sig_928 : std_logic;
	signal sig_929 : std_logic;
	signal sig_930 : std_logic;
	signal sig_931 : std_logic;
	signal sig_932 : std_logic;
	signal sig_933 : std_logic;
	signal sig_934 : std_logic;
	signal sig_935 : std_logic;
	signal sig_936 : std_logic;
	signal sig_937 : std_logic;
	signal sig_938 : std_logic;
	signal sig_939 : std_logic;
	signal sig_940 : std_logic;
	signal sig_941 : std_logic;
	signal sig_942 : std_logic;
	signal sig_943 : std_logic;
	signal sig_944 : std_logic;
	signal sig_945 : std_logic;
	signal sig_946 : std_logic;
	signal sig_947 : std_logic;
	signal sig_948 : std_logic;
	signal sig_949 : std_logic;
	signal sig_950 : std_logic;
	signal sig_951 : std_logic;
	signal sig_952 : std_logic;
	signal sig_953 : std_logic;
	signal sig_954 : std_logic;
	signal sig_955 : std_logic;
	signal sig_956 : std_logic;
	signal sig_957 : std_logic;
	signal sig_958 : std_logic;
	signal sig_959 : std_logic;
	signal sig_960 : std_logic;
	signal sig_961 : std_logic;
	signal sig_962 : std_logic;
	signal sig_963 : std_logic;
	signal sig_964 : std_logic;
	signal sig_965 : std_logic;
	signal sig_966 : std_logic;
	signal sig_967 : std_logic;
	signal sig_968 : std_logic;
	signal sig_969 : std_logic;
	signal sig_970 : std_logic;
	signal sig_971 : std_logic;
	signal sig_972 : std_logic;
	signal sig_973 : std_logic;
	signal sig_974 : std_logic;
	signal sig_975 : std_logic;
	signal sig_976 : std_logic;
	signal sig_977 : std_logic;
	signal sig_978 : std_logic;
	signal sig_979 : std_logic;
	signal sig_980 : std_logic;
	signal sig_981 : std_logic;
	signal sig_982 : std_logic;
	signal sig_983 : std_logic;
	signal sig_984 : std_logic;
	signal sig_985 : std_logic;
	signal sig_986 : std_logic;
	signal sig_987 : std_logic;
	signal sig_988 : std_logic;
	signal sig_989 : std_logic;
	signal sig_990 : std_logic;
	signal sig_991 : std_logic;
	signal sig_992 : std_logic;
	signal sig_993 : std_logic;
	signal sig_994 : std_logic;
	signal sig_995 : std_logic;
	signal sig_996 : std_logic;
	signal sig_997 : std_logic;
	signal sig_998 : std_logic;
	signal sig_999 : std_logic;
	signal sig_1000 : std_logic;
	signal sig_1001 : std_logic;
	signal sig_1002 : std_logic;
	signal sig_1003 : std_logic;
	signal sig_1004 : std_logic;
	signal sig_1005 : std_logic;
	signal sig_1006 : std_logic;
	signal sig_1007 : std_logic;
	signal sig_1008 : std_logic;
	signal sig_1009 : std_logic;
	signal sig_1010 : std_logic;
	signal sig_1011 : std_logic;
	signal sig_1012 : std_logic;
	signal sig_1013 : std_logic;
	signal sig_1014 : std_logic;
	signal sig_1015 : std_logic;
	signal sig_1016 : std_logic;
	signal sig_1017 : std_logic;
	signal sig_1018 : std_logic;
	signal sig_1019 : std_logic;
	signal sig_1020 : std_logic;
	signal sig_1021 : std_logic;
	signal sig_1022 : std_logic;
	signal sig_1023 : std_logic;
	signal sig_1024 : std_logic;
	signal sig_1025 : std_logic;
	signal sig_1026 : std_logic;
	signal sig_1027 : std_logic;
	signal sig_1028 : std_logic;
	signal sig_1029 : std_logic;
	signal sig_1030 : std_logic;
	signal sig_1031 : std_logic;
	signal sig_1032 : std_logic;
	signal sig_1033 : std_logic;
	signal sig_1034 : std_logic;
	signal sig_1035 : std_logic;
	signal sig_1036 : std_logic;
	signal sig_1037 : std_logic;
	signal sig_1038 : std_logic;
	signal sig_1039 : std_logic;
	signal sig_1040 : std_logic;
	signal sig_1041 : std_logic;
	signal sig_1042 : std_logic;
	signal sig_1043 : std_logic;
	signal sig_1044 : std_logic;
	signal sig_1045 : std_logic;
	signal sig_1046 : std_logic;
	signal sig_1047 : std_logic;
	signal sig_1048 : std_logic;
	signal sig_1049 : std_logic;
	signal sig_1050 : std_logic;
	signal sig_1051 : std_logic;
	signal sig_1052 : std_logic;
	signal sig_1053 : std_logic;
	signal sig_1054 : std_logic;
	signal sig_1055 : std_logic;
	signal sig_1056 : std_logic;
	signal sig_1057 : std_logic;
	signal sig_1058 : std_logic;
	signal sig_1059 : std_logic;
	signal sig_1060 : std_logic;
	signal sig_1061 : std_logic;
	signal sig_1062 : std_logic;
	signal sig_1063 : std_logic;
	signal sig_1064 : std_logic;
	signal sig_1065 : std_logic;
	signal sig_1066 : std_logic;
	signal sig_1067 : std_logic;
	signal sig_1068 : std_logic;
	signal sig_1069 : std_logic;
	signal sig_1070 : std_logic;
	signal sig_1071 : std_logic;
	signal sig_1072 : std_logic;
	signal sig_1073 : std_logic;
	signal sig_1074 : std_logic;
	signal sig_1075 : std_logic;
	signal sig_1076 : std_logic;
	signal sig_1077 : std_logic;
	signal sig_1078 : std_logic;
	signal sig_1079 : std_logic;
	signal sig_1080 : std_logic;
	signal sig_1081 : std_logic;
	signal sig_1082 : std_logic;
	signal sig_1083 : std_logic;
	signal sig_1084 : std_logic;
	signal sig_1085 : std_logic;
	signal sig_1086 : std_logic;
	signal sig_1087 : std_logic;
	signal sig_1088 : std_logic;
	signal sig_1089 : std_logic;
	signal sig_1090 : std_logic;
	signal sig_1091 : std_logic;
	signal sig_1092 : std_logic;
	signal sig_1093 : std_logic;
	signal sig_1094 : std_logic;
	signal sig_1095 : std_logic;
	signal sig_1096 : std_logic;
	signal sig_1097 : std_logic;
	signal sig_1098 : std_logic;
	signal sig_1099 : std_logic;
	signal sig_1100 : std_logic;
	signal sig_1101 : std_logic;
	signal sig_1102 : std_logic;
	signal sig_1103 : std_logic;
	signal sig_1104 : std_logic;
	signal sig_1105 : std_logic;
	signal sig_1106 : std_logic;
	signal sig_1107 : std_logic;
	signal sig_1108 : std_logic;
	signal sig_1109 : std_logic;
	signal sig_1110 : std_logic;
	signal sig_1111 : std_logic;
	signal sig_1112 : std_logic;
	signal sig_1113 : std_logic;
	signal sig_1114 : std_logic;
	signal sig_1115 : std_logic;
	signal sig_1116 : std_logic;
	signal sig_1117 : std_logic;
	signal sig_1118 : std_logic;
	signal sig_1119 : std_logic;
	signal sig_1120 : std_logic;
	signal sig_1121 : std_logic;
	signal sig_1122 : std_logic;
	signal sig_1123 : std_logic;
	signal sig_1124 : std_logic;
	signal sig_1125 : std_logic;
	signal sig_1126 : std_logic;
	signal sig_1127 : std_logic;
	signal sig_1128 : std_logic;
	signal sig_1129 : std_logic;
	signal sig_1130 : std_logic;
	signal sig_1131 : std_logic;
	signal sig_1132 : std_logic;
	signal sig_1133 : std_logic;
	signal sig_1134 : std_logic;
	signal sig_1135 : std_logic;
	signal sig_1136 : std_logic;
	signal sig_1137 : std_logic;
	signal sig_1138 : std_logic;
	signal sig_1139 : std_logic;
	signal sig_1140 : std_logic;
	signal sig_1141 : std_logic;
	signal sig_1142 : std_logic;
	signal sig_1143 : std_logic;
	signal sig_1144 : std_logic;
	signal sig_1145 : std_logic;
	signal sig_1146 : std_logic;
	signal sig_1147 : std_logic;
	signal sig_1148 : std_logic;
	signal sig_1149 : std_logic;
	signal sig_1150 : std_logic;
	signal sig_1151 : std_logic;
	signal sig_1152 : std_logic;
	signal sig_1153 : std_logic;
	signal sig_1154 : std_logic;
	signal sig_1155 : std_logic;
	signal sig_1156 : std_logic;
	signal sig_1157 : std_logic;
	signal sig_1158 : std_logic;
	signal sig_1159 : std_logic;
	signal sig_1160 : std_logic;
	signal sig_1161 : std_logic;
	signal sig_1162 : std_logic;
	signal sig_1163 : std_logic;
	signal sig_1164 : std_logic;
	signal sig_1165 : std_logic;
	signal sig_1166 : std_logic;
	signal sig_1167 : std_logic;
	signal sig_1168 : std_logic;
	signal sig_1169 : std_logic;
	signal sig_1170 : std_logic;
	signal sig_1171 : std_logic;
	signal sig_1172 : std_logic;
	signal sig_1173 : std_logic;
	signal sig_1174 : std_logic;
	signal sig_1175 : std_logic;
	signal sig_1176 : std_logic;
	signal sig_1177 : std_logic;
	signal sig_1178 : std_logic;
	signal sig_1179 : std_logic;
	signal sig_1180 : std_logic;
	signal sig_1181 : std_logic;
	signal sig_1182 : std_logic;
	signal sig_1183 : std_logic;
	signal sig_1184 : std_logic;
	signal sig_1185 : std_logic;
	signal sig_1186 : std_logic;
	signal sig_1187 : std_logic;
	signal sig_1188 : std_logic;
	signal sig_1189 : std_logic;
	signal sig_1190 : std_logic;
	signal sig_1191 : std_logic;
	signal sig_1192 : std_logic;
	signal sig_1193 : std_logic;
	signal sig_1194 : std_logic;
	signal sig_1195 : std_logic;
	signal sig_1196 : std_logic;
	signal sig_1197 : std_logic;
	signal sig_1198 : std_logic;
	signal sig_1199 : std_logic;
	signal sig_1200 : std_logic;
	signal sig_1201 : std_logic;
	signal sig_1202 : std_logic;
	signal sig_1203 : std_logic;
	signal sig_1204 : std_logic;
	signal sig_1205 : std_logic;
	signal sig_1206 : std_logic;
	signal sig_1207 : std_logic;
	signal sig_1208 : std_logic;
	signal sig_1209 : std_logic;
	signal sig_1210 : std_logic;
	signal sig_1211 : std_logic;
	signal sig_1212 : std_logic;
	signal sig_1213 : std_logic;
	signal sig_1214 : std_logic;
	signal sig_1215 : std_logic;
	signal sig_1216 : std_logic;
	signal sig_1217 : std_logic;
	signal sig_1218 : std_logic;
	signal sig_1219 : std_logic;
	signal sig_1220 : std_logic;
	signal sig_1221 : std_logic;
	signal sig_1222 : std_logic;
	signal sig_1223 : std_logic;
	signal sig_1224 : std_logic;
	signal sig_1225 : std_logic;
	signal sig_1226 : std_logic;
	signal sig_1227 : std_logic;
	signal sig_1228 : std_logic;
	signal sig_1229 : std_logic;
	signal sig_1230 : std_logic;
	signal sig_1231 : std_logic;
	signal sig_1232 : std_logic;
	signal sig_1233 : std_logic;
	signal sig_1234 : std_logic;
	signal sig_1235 : std_logic;
	signal sig_1236 : std_logic;
	signal sig_1237 : std_logic;
	signal sig_1238 : std_logic;
	signal sig_1239 : std_logic;
	signal sig_1240 : std_logic;
	signal sig_1241 : std_logic;
	signal sig_1242 : std_logic;
	signal sig_1243 : std_logic;
	signal sig_1244 : std_logic;
	signal sig_1245 : std_logic;
	signal sig_1246 : std_logic;
	signal sig_1247 : std_logic;
	signal sig_1248 : std_logic;
	signal sig_1249 : std_logic;
	signal sig_1250 : std_logic;
	signal sig_1251 : std_logic;
	signal sig_1252 : std_logic;
	signal sig_1253 : std_logic;
	signal sig_1254 : std_logic;
	signal sig_1255 : std_logic;
	signal sig_1256 : std_logic;
	signal sig_1257 : std_logic;
	signal sig_1258 : std_logic;
	signal sig_1259 : std_logic;
	signal sig_1260 : std_logic;
	signal sig_1261 : std_logic;
	signal sig_1262 : std_logic;
	signal sig_1263 : std_logic;
	signal sig_1264 : std_logic;
	signal sig_1265 : std_logic;
	signal sig_1266 : std_logic;
	signal sig_1267 : std_logic;
	signal sig_1268 : std_logic;
	signal sig_1269 : std_logic;
	signal sig_1270 : std_logic;
	signal sig_1271 : std_logic;
	signal sig_1272 : std_logic;
	signal sig_1273 : std_logic;
	signal sig_1274 : std_logic;
	signal sig_1275 : std_logic;
	signal sig_1276 : std_logic;
	signal sig_1277 : std_logic;
	signal sig_1278 : std_logic;
	signal sig_1279 : std_logic;
	signal sig_1280 : std_logic;
	signal sig_1281 : std_logic_vector(63 downto 0);
	signal sig_1282 : std_logic;
	signal sig_1283 : std_logic;
	signal sig_1284 : std_logic;
	signal sig_1285 : std_logic_vector(63 downto 0);
	signal sig_1286 : std_logic_vector(31 downto 0);
	signal sig_1287 : std_logic_vector(63 downto 0);
	signal sig_1288 : std_logic_vector(63 downto 0);
	signal sig_1289 : std_logic_vector(63 downto 0);
	signal sig_1290 : std_logic_vector(63 downto 0);
	signal sig_1291 : std_logic_vector(63 downto 0);
	signal sig_1292 : std_logic_vector(63 downto 0);
	signal sig_1293 : std_logic_vector(31 downto 0);
	signal sig_1294 : std_logic_vector(31 downto 0);
	signal sig_1295 : std_logic_vector(31 downto 0);
	signal sig_1296 : std_logic_vector(31 downto 0);
	signal sig_1297 : std_logic_vector(31 downto 0);
	signal sig_1298 : std_logic_vector(63 downto 0);
	signal sig_1299 : std_logic;
	signal sig_1300 : std_logic;
	signal sig_1301 : std_logic;
	signal sig_1302 : std_logic_vector(63 downto 0);
	signal sig_1303 : std_logic_vector(63 downto 0);
	signal sig_1304 : std_logic_vector(63 downto 0);
	signal sig_1305 : std_logic;
	signal sig_1306 : std_logic;
	signal sig_1307 : std_logic_vector(63 downto 0);
	signal sig_1308 : std_logic_vector(31 downto 0);
	signal sig_1309 : std_logic_vector(31 downto 0);
	signal sig_1310 : std_logic_vector(31 downto 0);
	signal sig_1311 : std_logic_vector(31 downto 0);
	signal sig_1312 : std_logic_vector(31 downto 0);
	signal sig_1313 : std_logic_vector(31 downto 0);
	signal sig_1314 : std_logic_vector(31 downto 0);
	signal sig_1315 : std_logic_vector(31 downto 0);
	signal sig_1316 : std_logic_vector(31 downto 0);
	signal sig_1317 : std_logic;
	signal sig_1318 : std_logic_vector(63 downto 0);
	signal sig_1319 : std_logic_vector(63 downto 0);

	-- Other inlined components

	signal and_757 : std_logic_vector(31 downto 0);
	signal or_758 : std_logic_vector(31 downto 0);
	signal and_760 : std_logic_vector(31 downto 0);
	signal or_761 : std_logic_vector(7 downto 0);
	signal not_762 : std_logic;
	signal not_764 : std_logic;
	signal not_766 : std_logic;
	signal or_767 : std_logic_vector(7 downto 0);
	signal mux_490 : std_logic_vector(30 downto 0);
	signal and_744 : std_logic_vector(31 downto 0);
	signal not_746 : std_logic;
	signal or_747 : std_logic_vector(31 downto 0);
	signal and_748 : std_logic_vector(31 downto 0);
	signal not_751 : std_logic;
	signal or_752 : std_logic_vector(31 downto 0);
	signal and_753 : std_logic_vector(31 downto 0);
	signal or_755 : std_logic_vector(31 downto 0);
	signal tqmf_reg0 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg1 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg2 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg3 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg4 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg5 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg6 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg7 : std_logic_vector(31 downto 0) := (others => '0');
	signal read32_buf_0 : std_logic_vector(31 downto 0) := (others => '0');
	signal write32_val_1 : std_logic_vector(31 downto 0) := (others => '0');
	signal filtez_zl : std_logic_vector(63 downto 0) := (others => '0');
	signal upzero_wd3 : std_logic_vector(31 downto 0) := (others => '0');
	signal upzero_wd2 : std_logic_vector(31 downto 0) := (others => '0');
	signal xh : std_logic_vector(31 downto 0) := (others => '0');
	signal or_714 : std_logic_vector(31 downto 0);
	signal and_715 : std_logic_vector(31 downto 0);
	signal and_723 : std_logic_vector(31 downto 0);
	signal and_727 : std_logic_vector(31 downto 0);
	signal not_728 : std_logic;
	signal and_735 : std_logic_vector(31 downto 0);
	signal or_742 : std_logic_vector(31 downto 0);
	signal and_743 : std_logic_vector(31 downto 0);
	signal xl : std_logic_vector(31 downto 0) := (others => '0');
	signal xd : std_logic_vector(31 downto 0) := (others => '0');
	signal xs : std_logic_vector(31 downto 0) := (others => '0');
	signal el : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_484 : std_logic_vector(31 downto 0);
	signal mux_486 : std_logic_vector(31 downto 0);
	signal sl : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_488 : std_logic_vector(30 downto 0);
	signal szl : std_logic_vector(31 downto 0) := (others => '0');
	signal il : std_logic_vector(5 downto 0) := (others => '0');
	signal mux_480 : std_logic_vector(31 downto 0);
	signal mux_476 : std_logic_vector(31 downto 0);
	signal mux_472 : std_logic_vector(30 downto 0);
	signal mux_474 : std_logic_vector(30 downto 0);
	signal mux_470 : std_logic_vector(31 downto 0);
	signal mux_468 : std_logic_vector(31 downto 0);
	signal mux_460 : std_logic_vector(31 downto 0);
	signal mux_462 : std_logic_vector(31 downto 0);
	signal nbl : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_456 : std_logic_vector(63 downto 0);
	signal al2 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_458 : std_logic_vector(31 downto 0);
	signal al1 : std_logic_vector(31 downto 0) := (others => '0');
	signal plt2 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_448 : std_logic_vector(31 downto 0);
	signal plt1 : std_logic_vector(31 downto 0) := (others => '0');
	signal plt : std_logic_vector(31 downto 0) := (others => '0');
	signal dlt : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_434 : std_logic_vector(31 downto 0);
	signal rlt2 : std_logic_vector(30 downto 0) := (others => '0');
	signal mux_438 : std_logic_vector(31 downto 0);
	signal rlt1 : std_logic_vector(30 downto 0) := (others => '0');
	signal mux_440 : std_logic_vector(31 downto 0);
	signal rlt : std_logic_vector(30 downto 0) := (others => '0');
	signal mux_430 : std_logic_vector(31 downto 0);
	signal mux_432 : std_logic_vector(31 downto 0);
	signal detl : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_424 : std_logic_vector(31 downto 0);
	signal mux_426 : std_logic_vector(31 downto 0);
	signal mux_422 : std_logic_vector(31 downto 0);
	signal deth : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_416 : std_logic_vector(63 downto 0);
	signal sh : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_414 : std_logic_vector(63 downto 0);
	signal eh : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_406 : std_logic_vector(63 downto 0);
	signal mux_400 : std_logic_vector(31 downto 0);
	signal mux_402 : std_logic_vector(63 downto 0);
	signal ih : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_403 : std_logic_vector(63 downto 0);
	signal mux_404 : std_logic_vector(63 downto 0);
	signal dh : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_395 : std_logic_vector(63 downto 0);
	signal mux_396 : std_logic_vector(63 downto 0);
	signal mux_397 : std_logic_vector(63 downto 0);
	signal mux_398 : std_logic_vector(31 downto 0);
	signal mux_399 : std_logic_vector(63 downto 0);
	signal nbh : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_383 : std_logic_vector(5 downto 0);
	signal rh : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_385 : std_logic_vector(6 downto 0);
	signal yh : std_logic_vector(30 downto 0) := (others => '0');
	signal mux_390 : std_logic_vector(63 downto 0);
	signal ph : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_391 : std_logic_vector(63 downto 0);
	signal mux_376 : std_logic_vector(6 downto 0);
	signal mux_377 : std_logic_vector(31 downto 0);
	signal mux_372 : std_logic_vector(31 downto 0);
	signal ah2 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_374 : std_logic_vector(6 downto 0);
	signal ah1 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_364 : std_logic_vector(31 downto 0);
	signal mux_365 : std_logic_vector(32 downto 0);
	signal mux_366 : std_logic_vector(31 downto 0);
	signal ph2 : std_logic_vector(31 downto 0) := (others => '0');
	signal ph1 : std_logic_vector(31 downto 0) := (others => '0');
	signal rh2 : std_logic_vector(30 downto 0) := (others => '0');
	signal mux_363 : std_logic_vector(32 downto 0);
	signal rh1 : std_logic_vector(30 downto 0) := (others => '0');
	signal mux_352 : std_logic_vector(63 downto 0);
	signal mux_353 : std_logic_vector(63 downto 0);
	signal mux_354 : std_logic_vector(63 downto 0);
	signal rl : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_355 : std_logic_vector(63 downto 0);
	signal mux_356 : std_logic_vector(63 downto 0);
	signal dec_dlt : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_detl : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_349 : std_logic_vector(32 downto 0);
	signal mux_350 : std_logic_vector(31 downto 0);
	signal mux_351 : std_logic_vector(63 downto 0);
	signal dec_deth : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_341 : std_logic_vector(63 downto 0);
	signal mux_342 : std_logic_vector(63 downto 0);
	signal mux_338 : std_logic_vector(31 downto 0);
	signal dec_plt2 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_plt1 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_336 : std_logic_vector(31 downto 0);
	signal dec_plt : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_320 : std_logic_vector(31 downto 0);
	signal dec_sl : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_322 : std_logic_vector(31 downto 0);
	signal mux_324 : std_logic_vector(31 downto 0);
	signal mux_326 : std_logic_vector(31 downto 0);
	signal mux_310 : std_logic_vector(31 downto 0);
	signal dec_rlt : std_logic_vector(30 downto 0) := (others => '0');
	signal mux_314 : std_logic_vector(32 downto 0);
	signal mux_315 : std_logic_vector(31 downto 0);
	signal dec_rlt2 : std_logic_vector(30 downto 0) := (others => '0');
	signal mux_316 : std_logic_vector(31 downto 0);
	signal mux_318 : std_logic_vector(31 downto 0);
	signal dec_rlt1 : std_logic_vector(30 downto 0) := (others => '0');
	signal dec_al2 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_308 : std_logic_vector(31 downto 0);
	signal dec_al1 : std_logic_vector(31 downto 0) := (others => '0');
	signal dl : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_292 : std_logic_vector(31 downto 0);
	signal mux_294 : std_logic_vector(31 downto 0);
	signal dec_nbh : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_296 : std_logic_vector(31 downto 0);
	signal dec_dh : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_298 : std_logic_vector(31 downto 0);
	signal dec_nbl : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_290 : std_logic_vector(31 downto 0);
	signal mux_286 : std_logic_vector(31 downto 0);
	signal mux_288 : std_logic_vector(31 downto 0);
	signal mux_284 : std_logic_vector(31 downto 0);
	signal mux_278 : std_logic_vector(31 downto 0);
	signal dec_rh2 : std_logic_vector(30 downto 0) := (others => '0');
	signal mux_280 : std_logic_vector(31 downto 0);
	signal mux_282 : std_logic_vector(31 downto 0);
	signal dec_rh1 : std_logic_vector(30 downto 0) := (others => '0');
	signal mux_272 : std_logic_vector(31 downto 0);
	signal dec_ah2 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_274 : std_logic_vector(31 downto 0);
	signal mux_276 : std_logic_vector(31 downto 0);
	signal dec_ah1 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_ph : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_262 : std_logic_vector(31 downto 0);
	signal dec_sh : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_ph2 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_260 : std_logic_vector(31 downto 0);
	signal dec_ph1 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_250 : std_logic_vector(31 downto 0);
	signal abs_m_3 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_248 : std_logic_vector(31 downto 0);
	signal mux_244 : std_logic_vector(31 downto 0);
	signal mux_246 : std_logic_vector(31 downto 0);
	signal mux_242 : std_logic_vector(31 downto 0);
	signal mux_238 : std_logic_vector(31 downto 0);
	signal mux_240 : std_logic_vector(31 downto 0);
	signal filtep_pl_14 : std_logic_vector(63 downto 0) := (others => '0');
	signal mux_236 : std_logic_vector(31 downto 0);
	signal quantl_el_16 : std_logic := '0';
	signal mux_232 : std_logic_vector(31 downto 0);
	signal mux_234 : std_logic_vector(31 downto 0);
	signal quantl_detl_17 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_230 : std_logic_vector(31 downto 0);
	signal quantl_ril_18 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_226 : std_logic_vector(31 downto 0);
	signal mux_228 : std_logic_vector(31 downto 0);
	signal quantl_mil_19 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_224 : std_logic_vector(31 downto 0);
	signal quantl_wd_20 : std_logic_vector(63 downto 0) := (others => '0');
	signal mux_220 : std_logic_vector(31 downto 0);
	signal mux_222 : std_logic_vector(31 downto 0);
	signal quantl_decis_21 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_218 : std_logic_vector(31 downto 0);
	signal logscl_nbl_27 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_214 : std_logic_vector(31 downto 0);
	signal mux_216 : std_logic_vector(31 downto 0);
	signal logscl_wd_28 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_212 : std_logic_vector(31 downto 0);
	signal mux_208 : std_logic_vector(31 downto 0);
	signal mux_210 : std_logic_vector(31 downto 0);
	signal mux_206 : std_logic_vector(31 downto 0);
	signal mux_202 : std_logic_vector(31 downto 0);
	signal mux_204 : std_logic_vector(31 downto 0);
	signal scalel_wd3_35 : std_logic_vector(28 downto 0) := (others => '0');
	signal mux_200 : std_logic_vector(31 downto 0);
	signal mux_196 : std_logic_vector(31 downto 0);
	signal mux_198 : std_logic_vector(31 downto 0);
	signal mux_194 : std_logic_vector(31 downto 0);
	signal mux_190 : std_logic_vector(31 downto 0);
	signal mux_192 : std_logic_vector(31 downto 0);
	signal mux_188 : std_logic_vector(31 downto 0);
	signal mux_184 : std_logic_vector(31 downto 0);
	signal mux_186 : std_logic_vector(31 downto 0);
	signal uppol2_wd4_42 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_182 : std_logic_vector(31 downto 0);
	signal uppol2_apl2_43 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_178 : std_logic_vector(31 downto 0);
	signal mux_180 : std_logic_vector(31 downto 0);
	signal mux_176 : std_logic_vector(31 downto 0);
	signal mux_172 : std_logic_vector(31 downto 0);
	signal mux_174 : std_logic_vector(31 downto 0);
	signal mux_170 : std_logic_vector(31 downto 0);
	signal uppol1_wd2_51 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_166 : std_logic_vector(31 downto 0);
	signal mux_168 : std_logic_vector(31 downto 0);
	signal uppol1_wd3_52 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_164 : std_logic_vector(31 downto 0);
	signal uppol1_apl1_53 : std_logic_vector(31 downto 0) := (others => '0');
	signal logsch_nbh_57 : std_logic_vector(31 downto 0) := (others => '0');
	signal logsch_wd_58 : std_logic_vector(31 downto 0) := (others => '0');
	signal encode_xin1_61 : std_logic_vector(31 downto 0) := (others => '0');
	signal encode_xin2_62 : std_logic_vector(31 downto 0) := (others => '0');
	signal encode_xa_67 : std_logic_vector(63 downto 0) := (others => '0');
	signal encode_xb_68 : std_logic_vector(63 downto 0) := (others => '0');
	signal encode_decis_69 : std_logic_vector(31 downto 0) := (others => '0');
	signal not_709 : std_logic;
	signal or_710 : std_logic_vector(31 downto 0);
	signal decode_input_98 : std_logic_vector(29 downto 0) := (others => '0');
	signal decode_xa1_100 : std_logic_vector(63 downto 0) := (others => '0');
	signal decode_xa2_101 : std_logic_vector(63 downto 0) := (others => '0');
	signal or_692 : std_logic_vector(7 downto 0);
	signal not_693 : std_logic;
	signal augh_main_i_132 : std_logic_vector(31 downto 0) := (others => '0');
	signal encode_ret0_136 : std_logic_vector(31 downto 0) := (others => '0');
	signal not_768 : std_logic;
	signal or_769 : std_logic_vector(31 downto 0);
	signal and_770 : std_logic_vector(31 downto 0);
	signal and_771 : std_logic_vector(31 downto 0);
	signal or_619 : std_logic_vector(7 downto 0);
	signal not_620 : std_logic;
	signal or_621 : std_logic_vector(7 downto 0);
	signal not_622 : std_logic;
	signal or_623 : std_logic_vector(7 downto 0);
	signal not_624 : std_logic;
	signal or_625 : std_logic_vector(7 downto 0);
	signal not_626 : std_logic;
	signal or_627 : std_logic_vector(7 downto 0);
	signal and_633 : std_logic_vector(31 downto 0);
	signal not_628 : std_logic;
	signal or_629 : std_logic_vector(7 downto 0);
	signal not_630 : std_logic;
	signal dec_del_dhx_reg0 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_dhx_reg1 : std_logic_vector(31 downto 0) := (others => '0');
	signal or_631 : std_logic_vector(31 downto 0);
	signal or_634 : std_logic_vector(7 downto 0);
	signal not_635 : std_logic;
	signal or_636 : std_logic_vector(7 downto 0);
	signal not_637 : std_logic;
	signal dec_del_bph_reg0 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_bph_reg1 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_bph_reg2 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_bph_reg3 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_bph_reg4 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_bph_reg5 : std_logic_vector(31 downto 0) := (others => '0');
	signal and_632 : std_logic_vector(31 downto 0);
	signal or_641 : std_logic_vector(31 downto 0);
	signal and_640 : std_logic_vector(31 downto 0);
	signal and_645 : std_logic_vector(31 downto 0);
	signal and_639 : std_logic_vector(31 downto 0);
	signal and_643 : std_logic_vector(31 downto 0);
	signal and_650 : std_logic_vector(31 downto 0);
	signal or_651 : std_logic_vector(31 downto 0);
	signal or_644 : std_logic_vector(31 downto 0);
	signal and_649 : std_logic_vector(31 downto 0);
	signal dec_del_dltx_reg0 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_dltx_reg1 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_498 : std_logic_vector(31 downto 0);
	signal mux_500 : std_logic_vector(31 downto 0);
	signal mux_502 : std_logic_vector(31 downto 0);
	signal mux_504 : std_logic_vector(31 downto 0);
	signal and_652 : std_logic_vector(31 downto 0);
	signal and_653 : std_logic_vector(31 downto 0);
	signal or_654 : std_logic_vector(31 downto 0);
	signal and_655 : std_logic_vector(31 downto 0);
	signal and_656 : std_logic_vector(31 downto 0);
	signal or_657 : std_logic_vector(31 downto 0);
	signal and_658 : std_logic_vector(31 downto 0);
	signal and_659 : std_logic_vector(31 downto 0);
	signal dec_del_bpl_reg0 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_bpl_reg1 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_bpl_reg2 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_bpl_reg3 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_bpl_reg4 : std_logic_vector(31 downto 0) := (others => '0');
	signal dec_del_bpl_reg5 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_510 : std_logic_vector(30 downto 0);
	signal mux_512 : std_logic_vector(30 downto 0);
	signal not_661 : std_logic;
	signal and_665 : std_logic_vector(31 downto 0);
	signal or_666 : std_logic_vector(31 downto 0);
	signal delay_bph_reg0 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_bph_reg1 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_bph_reg2 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_bph_reg3 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_bph_reg4 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_bph_reg5 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_514 : std_logic_vector(31 downto 0);
	signal mux_516 : std_logic_vector(31 downto 0);
	signal mux_518 : std_logic_vector(31 downto 0);
	signal mux_520 : std_logic_vector(31 downto 0);
	signal and_647 : std_logic_vector(31 downto 0);
	signal and_664 : std_logic_vector(31 downto 0);
	signal and_667 : std_logic_vector(31 downto 0);
	signal and_670 : std_logic_vector(31 downto 0);
	signal and_672 : std_logic_vector(31 downto 0);
	signal or_674 : std_logic_vector(31 downto 0);
	signal delay_dhx_reg0 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_dhx_reg1 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_528 : std_logic_vector(31 downto 0);
	signal or_638 : std_logic_vector(31 downto 0);
	signal and_642 : std_logic_vector(31 downto 0);
	signal or_648 : std_logic_vector(31 downto 0);
	signal or_669 : std_logic_vector(31 downto 0);
	signal and_676 : std_logic_vector(31 downto 0);
	signal delay_dltx_reg0 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_dltx_reg1 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_532 : std_logic_vector(31 downto 0);
	signal mux_534 : std_logic_vector(1 downto 0);
	signal mux_535 : std_logic_vector(1 downto 0);
	signal or_663 : std_logic_vector(31 downto 0);
	signal and_668 : std_logic_vector(31 downto 0);
	signal or_679 : std_logic_vector(7 downto 0);
	signal not_680 : std_logic;
	signal not_682 : std_logic;
	signal or_683 : std_logic_vector(7 downto 0);
	signal and_686 : std_logic_vector(31 downto 0);
	signal and_689 : std_logic_vector(31 downto 0);
	signal delay_bpl_reg0 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_bpl_reg1 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_bpl_reg2 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_bpl_reg3 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_bpl_reg4 : std_logic_vector(31 downto 0) := (others => '0');
	signal delay_bpl_reg5 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_540 : std_logic_vector(31 downto 0);
	signal mux_544 : std_logic_vector(31 downto 0);
	signal or_660 : std_logic_vector(7 downto 0);
	signal or_677 : std_logic_vector(7 downto 0);
	signal not_678 : std_logic;
	signal not_684 : std_logic;
	signal or_685 : std_logic_vector(31 downto 0);
	signal or_688 : std_logic_vector(31 downto 0);
	signal or_695 : std_logic_vector(7 downto 0);
	signal accumc_reg0 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumc_reg1 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumc_reg2 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumc_reg3 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumc_reg4 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumc_reg5 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumc_reg6 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumc_reg7 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumc_reg8 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumc_reg9 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumc_reg10 : std_logic_vector(31 downto 0) := (others => '0');
	signal not_671 : std_logic;
	signal not_696 : std_logic;
	signal or_697 : std_logic_vector(7 downto 0);
	signal not_698 : std_logic;
	signal or_699 : std_logic_vector(25 downto 0);
	signal not_703 : std_logic;
	signal accumd_reg0 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumd_reg1 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumd_reg2 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumd_reg3 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumd_reg4 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumd_reg5 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumd_reg6 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumd_reg7 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumd_reg8 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumd_reg9 : std_logic_vector(31 downto 0) := (others => '0');
	signal accumd_reg10 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_563 : std_logic_vector(31 downto 0);
	signal mux_549 : std_logic_vector(30 downto 0);
	signal mux_551 : std_logic_vector(30 downto 0);
	signal mux_557 : std_logic_vector(31 downto 0);
	signal mux_559 : std_logic_vector(31 downto 0);
	signal mux_561 : std_logic_vector(31 downto 0);
	signal not_646 : std_logic;
	signal and_675 : std_logic_vector(31 downto 0);
	signal and_681 : std_logic_vector(31 downto 0);
	signal not_690 : std_logic;
	signal and_691 : std_logic_vector(31 downto 0);
	signal and_702 : std_logic_vector(31 downto 0);
	signal or_705 : std_logic_vector(31 downto 0);
	signal not_712 : std_logic;
	signal or_717 : std_logic_vector(31 downto 0);
	signal not_722 : std_logic;
	signal tqmf_reg8 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg9 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg10 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg11 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg12 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg13 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg14 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg15 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg16 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg17 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg18 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg19 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg20 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg21 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_565 : std_logic_vector(31 downto 0);
	signal mux_567 : std_logic_vector(4 downto 0);
	signal mux_568 : std_logic_vector(3 downto 0);
	signal mux_570 : std_logic_vector(3 downto 0);
	signal and_687 : std_logic_vector(31 downto 0);
	signal and_704 : std_logic_vector(31 downto 0);
	signal and_707 : std_logic_vector(31 downto 0);
	signal and_716 : std_logic_vector(31 downto 0);
	signal or_720 : std_logic_vector(31 downto 0);
	signal and_721 : std_logic_vector(31 downto 0);
	signal and_724 : std_logic_vector(31 downto 0);
	signal or_730 : std_logic_vector(7 downto 0);
	signal not_731 : std_logic;
	signal or_732 : std_logic_vector(7 downto 0);
	signal not_733 : std_logic;
	signal or_734 : std_logic_vector(31 downto 0);
	signal or_740 : std_logic_vector(7 downto 0);
	signal not_741 : std_logic;
	signal and_706 : std_logic_vector(31 downto 0);
	signal and_713 : std_logic_vector(31 downto 0);
	signal and_718 : std_logic_vector(31 downto 0);
	signal and_719 : std_logic_vector(31 downto 0);
	signal not_725 : std_logic;
	signal or_726 : std_logic_vector(31 downto 0);
	signal tqmf_reg22 : std_logic_vector(31 downto 0) := (others => '0');
	signal tqmf_reg23 : std_logic_vector(31 downto 0) := (others => '0');
	signal mux_587 : std_logic_vector(31 downto 0);
	signal mux_589 : std_logic_vector(31 downto 0);
	signal mux_591 : std_logic_vector(63 downto 0);
	signal mux_593 : std_logic_vector(31 downto 0);
	signal mux_597 : std_logic_vector(31 downto 0);
	signal mux_599 : std_logic_vector(31 downto 0);
	signal mux_601 : std_logic_vector(31 downto 0);
	signal mux_603 : std_logic_vector(31 downto 0);
	signal mux_605 : std_logic_vector(31 downto 0);
	signal mux_607 : std_logic_vector(31 downto 0);
	signal mux_609 : std_logic_vector(31 downto 0);
	signal mux_611 : std_logic_vector(31 downto 0);
	signal or_701 : std_logic_vector(31 downto 0);
	signal or_708 : std_logic_vector(7 downto 0);
	signal and_711 : std_logic_vector(31 downto 0);
	signal and_729 : std_logic_vector(31 downto 0);
	signal and_736 : std_logic_vector(31 downto 0);
	signal or_737 : std_logic_vector(31 downto 0);
	signal and_738 : std_logic_vector(31 downto 0);
	signal and_739 : std_logic_vector(31 downto 0);
	signal or_745 : std_logic_vector(7 downto 0);
	signal and_749 : std_logic_vector(31 downto 0);
	signal and_750 : std_logic_vector(31 downto 0);
	signal and_754 : std_logic_vector(31 downto 0);
	signal and_756 : std_logic_vector(31 downto 0);
	signal and_759 : std_logic_vector(31 downto 0);
	signal and_763 : std_logic_vector(31 downto 0);
	signal or_765 : std_logic_vector(7 downto 0);
	signal or_772 : std_logic_vector(7 downto 0);
	signal not_773 : std_logic;
	signal or_774 : std_logic_vector(7 downto 0);
	signal not_775 : std_logic;
	signal or_776 : std_logic_vector(7 downto 0);
	signal not_777 : std_logic;
	signal or_778 : std_logic_vector(7 downto 0);
	signal not_779 : std_logic;
	signal or_780 : std_logic_vector(7 downto 0);
	signal not_781 : std_logic;

	-- This utility function is used for inlining MUX behaviour

	-- Little utility function to ease concatenation of an std_logic
	-- and explicitely return an std_logic_vector
	function repeat(N: natural; B: std_logic) return std_logic_vector is
		variable result: std_logic_vector(N-1 downto 0);
	begin
		result := (others => B);
		return result;
	end;

begin

	-- Instantiation of components

	sub_147_i : sub_147 port map (
		output => sig_1318,
		sign => '1',
		ge => sig_1317,
		in_a => sig_1319,
		in_b => "1111111111111111111111111111111111111111111111111101000000000000"
	);

	qq4_code4_table_i : qq4_code4_table port map (
		clk => sig_clock,
		ra0_data => sig_1316,
		ra0_addr => mux_570
	);

	qq6_code6_table_i : qq6_code6_table port map (
		clk => sig_clock,
		ra0_data => sig_1315,
		ra0_addr => il
	);

	wl_code_table_i : wl_code_table port map (
		clk => sig_clock,
		ra0_data => sig_1314,
		ra0_addr => mux_568
	);

	ilb_table_i : ilb_table port map (
		clk => sig_clock,
		ra0_data => sig_1313,
		ra0_addr => mux_567
	);

	decis_levl_i : decis_levl port map (
		clk => sig_clock,
		ra0_data => sig_1312,
		ra0_addr => quantl_mil_19(4 downto 0)
	);

	quant26bt_pos_i : quant26bt_pos port map (
		clk => sig_clock,
		ra0_data => sig_1311,
		ra0_addr => quantl_mil_19(4 downto 0)
	);

	quant26bt_neg_i : quant26bt_neg port map (
		clk => sig_clock,
		ra0_data => sig_1310,
		ra0_addr => quantl_mil_19(4 downto 0)
	);

	qq2_code2_table_i : qq2_code2_table port map (
		clk => sig_clock,
		ra0_data => sig_1309,
		ra0_addr => mux_535
	);

	wh_code_table_i : wh_code_table port map (
		clk => sig_clock,
		ra0_data => sig_1308,
		ra0_addr => mux_534
	);

	cmp_694_i : cmp_694 port map (
		in1 => dlt,
		in0 => "00000000000000000000000000000000",
		eq => augh_test_78
	);

	cmp_700_i : cmp_700 port map (
		in1 => dec_dh,
		in0 => "00000000000000000000000000000000",
		eq => augh_test_124
	);

	sub_144_i : sub_144 port map (
		output => sig_1307,
		le => sig_1306,
		sign => '1',
		ge => sig_1305,
		in_a => mux_402,
		in_b => mux_403
	);

	mul_145_i : mul_145 port map (
		output => sig_1304,
		in_a => mux_399,
		in_b => mux_400
	);

	mul_146_i : mul_146 port map (
		output => sig_1303,
		in_a => mux_397,
		in_b => mux_398
	);

	sub_143_i : sub_143 port map (
		output => sig_1302,
		lt => sig_1301,
		le => sig_1300,
		sign => '1',
		gt => sig_1299,
		in_a => mux_395,
		in_b => mux_396
	);

	add_142_i : add_142 port map (
		output => sig_1298,
		in_a => mux_390,
		in_b => mux_391
	);

	test_data_i : test_data port map (
		clk => sig_clock,
		ra0_data => sig_1297,
		wa0_addr => mux_385,
		wa0_en => sig_1213,
		ra0_addr => sig_1298(6 downto 0),
		wa0_data => read32_buf_0,
		ra1_data => sig_1296,
		ra1_addr => augh_main_i_132(6 downto 0)
	);

	shr_141_i : shr_141 port map (
		output => sig_1295,
		input => sig_1313,
		shift => mux_383,
		padding => sig_1313(31)
	);

	compressed_i : compressed port map (
		clk => sig_clock,
		ra0_data => sig_1294,
		wa0_addr => augh_main_i_132(7 downto 1),
		wa0_en => sig_1020,
		ra0_addr => augh_main_i_132(7 downto 1),
		wa0_data => encode_ret0_136
	);

	result_i : result port map (
		clk => sig_clock,
		ra0_data => sig_1293,
		wa0_addr => mux_374,
		wa0_en => sig_1088,
		ra0_addr => mux_376,
		wa0_data => mux_377
	);

	cmp_662_i : cmp_662 port map (
		in1 => dec_dlt,
		in0 => "00000000000000000000000000000000",
		eq => augh_test_113
	);

	cmp_673_i : cmp_673 port map (
		in1 => dh,
		in0 => "00000000000000000000000000000000",
		eq => augh_test_92
	);

	mul_148_i : mul_148 port map (
		output => sig_1292,
		in_a => mux_365,
		in_b => mux_366
	);

	mul_149_i : mul_149 port map (
		output => sig_1291,
		in_a => mux_363,
		in_b => mux_364
	);

	add_153_i : add_153 port map (
		output => sig_1290,
		in_a => mux_355,
		in_b => mux_356
	);

	add_154_i : add_154 port map (
		output => sig_1289,
		in_a => mux_353,
		in_b => mux_354
	);

	add_155_i : add_155 port map (
		output => sig_1288,
		in_a => mux_351,
		in_b => mux_352
	);

	mul_156_i : mul_156 port map (
		output => sig_1287,
		in_a => mux_349,
		in_b => mux_350
	);

	add_159_i : add_159 port map (
		output => sig_1286,
		in_a => uppol2_wd4_42,
		in_b => sig_1281(38 downto 7)
	);

	sub_160_i : sub_160 port map (
		output => sig_1285,
		lt => sig_1284,
		le => sig_1283,
		sign => '1',
		ge => sig_1282,
		in_a => mux_341,
		in_b => mux_342
	);

	mul_161_i : mul_161 port map (
		output => sig_1281,
		in_a => mux_314,
		in_b => mux_315
	);

	fsm_163_i : fsm_163 port map (
		clock => sig_clock,
		reset => sig_reset,
		out91 => sig_1280,
		out92 => sig_1279,
		out93 => sig_1278,
		in7 => augh_test_138,
		out94 => sig_1277,
		out95 => sig_1276,
		out98 => sig_1275,
		out100 => sig_1274,
		out101 => sig_1273,
		out102 => sig_1272,
		out104 => sig_1271,
		out105 => sig_1270,
		out106 => sig_1269,
		out107 => sig_1268,
		out108 => sig_1267,
		out109 => sig_1266,
		out111 => sig_1265,
		out114 => sig_1264,
		out116 => sig_1263,
		out118 => sig_1262,
		out119 => sig_1261,
		out120 => sig_1260,
		out128 => sig_1259,
		out130 => sig_1258,
		out131 => sig_1257,
		out132 => sig_1256,
		out137 => sig_1255,
		in8 => augh_test_137,
		out152 => sig_1254,
		out155 => sig_1253,
		out156 => sig_1252,
		out31 => sig_1251,
		in2 => sig_start,
		out28 => sig_1250,
		out29 => sig_1249,
		out30 => sig_1248,
		out26 => sig_1247,
		out27 => sig_1246,
		out24 => sig_1245,
		out25 => sig_1244,
		out77 => sig_1243,
		out79 => sig_1242,
		out80 => sig_1241,
		out82 => sig_1240,
		out34 => sig_1239,
		out35 => sig_1238,
		out36 => sig_1237,
		out32 => sig_1236,
		out33 => sig_1235,
		out40 => sig_1234,
		out41 => sig_1233,
		out88 => sig_1232,
		out89 => sig_1231,
		out21 => sig_1230,
		out22 => sig_1229,
		out23 => sig_1228,
		out73 => sig_1227,
		out76 => sig_1226,
		in6 => augh_test_124,
		out70 => sig_1225,
		out12 => sig_1224,
		out13 => sig_1223,
		out14 => sig_1222,
		out17 => sig_1221,
		out18 => sig_1220,
		out19 => sig_1219,
		out20 => sig_1218,
		out9 => sig_1217,
		out11 => stdout_rdy,
		out8 => sig_1216,
		out2 => sig_1215,
		out4 => sig_1214,
		out5 => sig_1213,
		in1 => stdin_ack,
		out6 => sig_1212,
		out7 => sig_1211,
		out0 => sig_1210,
		out1 => sig_1209,
		out37 => sig_1208,
		out38 => sig_1207,
		out39 => sig_1206,
		out1222 => sig_1205,
		out1223 => sig_1204,
		out1224 => sig_1203,
		out1225 => sig_1202,
		out1226 => sig_1201,
		out1228 => sig_1200,
		out1230 => sig_1199,
		in0 => stdout_ack,
		out67 => sig_1198,
		out68 => sig_1197,
		out65 => sig_1196,
		out66 => sig_1195,
		in5 => augh_test_78,
		out62 => sig_1194,
		out58 => sig_1193,
		out56 => sig_1192,
		in4 => augh_test_92,
		out57 => sig_1191,
		out54 => sig_1190,
		out55 => sig_1189,
		out51 => sig_1188,
		out52 => sig_1187,
		out53 => sig_1186,
		in3 => augh_test_113,
		out46 => sig_1185,
		out47 => sig_1184,
		out48 => sig_1183,
		out49 => sig_1182,
		out50 => sig_1181,
		out42 => sig_1180,
		out43 => sig_1179,
		out44 => sig_1178,
		out45 => sig_1177,
		in9 => augh_test_23,
		in10 => augh_test_24,
		out171 => sig_1176,
		in11 => augh_test_135,
		out191 => sig_1175,
		out207 => sig_1174,
		out208 => sig_1173,
		out209 => sig_1172,
		out212 => sig_1171,
		out213 => sig_1170,
		out216 => sig_1169,
		out220 => sig_1168,
		out221 => sig_1167,
		out223 => sig_1166,
		out224 => sig_1165,
		out226 => sig_1164,
		out227 => sig_1163,
		out228 => sig_1162,
		out229 => sig_1161,
		out230 => sig_1160,
		out233 => sig_1159,
		out235 => sig_1158,
		out236 => sig_1157,
		out237 => sig_1156,
		out238 => sig_1155,
		out239 => sig_1154,
		out241 => sig_1153,
		out250 => sig_1152,
		out258 => sig_1151,
		out259 => sig_1150,
		out261 => sig_1149,
		out270 => sig_1148,
		out276 => sig_1147,
		out277 => sig_1146,
		out283 => sig_1145,
		out285 => sig_1144,
		out287 => sig_1143,
		out290 => sig_1142,
		out291 => sig_1141,
		out293 => sig_1140,
		out301 => sig_1139,
		out303 => sig_1138,
		out304 => sig_1137,
		out315 => sig_1136,
		out319 => sig_1135,
		out321 => sig_1134,
		out330 => sig_1133,
		out335 => sig_1132,
		out338 => sig_1131,
		out341 => sig_1130,
		out342 => sig_1129,
		out344 => sig_1128,
		out347 => sig_1127,
		out351 => sig_1126,
		out354 => sig_1125,
		out355 => sig_1124,
		out356 => sig_1123,
		out357 => sig_1122,
		out358 => sig_1121,
		out360 => sig_1120,
		out361 => sig_1119,
		out362 => sig_1118,
		out365 => sig_1117,
		out367 => sig_1116,
		out368 => sig_1115,
		out370 => sig_1114,
		out375 => sig_1113,
		out376 => sig_1112,
		out378 => sig_1111,
		out381 => sig_1110,
		out382 => sig_1109,
		out386 => sig_1108,
		out387 => sig_1107,
		out388 => sig_1106,
		out390 => sig_1105,
		out392 => sig_1104,
		out393 => sig_1103,
		out394 => sig_1102,
		out397 => sig_1101,
		out403 => sig_1100,
		out404 => sig_1099,
		out408 => sig_1098,
		out409 => sig_1097,
		out410 => sig_1096,
		out412 => sig_1095,
		out416 => sig_1094,
		out417 => sig_1093,
		out418 => sig_1092,
		out419 => sig_1091,
		out420 => sig_1090,
		out421 => sig_1089,
		out424 => sig_1088,
		out425 => sig_1087,
		out430 => sig_1086,
		out431 => sig_1085,
		out434 => sig_1084,
		out436 => sig_1083,
		out438 => sig_1082,
		out439 => sig_1081,
		out440 => sig_1080,
		out441 => sig_1079,
		out442 => sig_1078,
		out443 => sig_1077,
		out444 => sig_1076,
		out445 => sig_1075,
		out446 => sig_1074,
		out447 => sig_1073,
		out448 => sig_1072,
		out450 => sig_1071,
		out451 => sig_1070,
		out454 => sig_1069,
		out457 => sig_1068,
		out460 => sig_1067,
		out463 => sig_1066,
		out465 => sig_1065,
		out466 => sig_1064,
		out472 => sig_1063,
		out473 => sig_1062,
		out475 => sig_1061,
		out476 => sig_1060,
		out479 => sig_1059,
		out480 => sig_1058,
		out481 => sig_1057,
		out482 => sig_1056,
		out484 => sig_1055,
		out485 => sig_1054,
		out489 => sig_1053,
		out491 => sig_1052,
		out494 => sig_1051,
		out497 => sig_1050,
		out500 => sig_1049,
		out503 => sig_1048,
		out504 => sig_1047,
		out505 => sig_1046,
		out508 => sig_1045,
		out509 => sig_1044,
		out513 => sig_1043,
		out514 => sig_1042,
		out516 => sig_1041,
		out521 => sig_1040,
		out523 => sig_1039,
		out524 => sig_1038,
		out525 => sig_1037,
		out530 => sig_1036,
		out532 => sig_1035,
		out533 => sig_1034,
		out535 => sig_1033,
		out536 => sig_1032,
		out539 => sig_1031,
		out541 => sig_1030,
		out543 => sig_1029,
		out545 => sig_1028,
		out547 => sig_1027,
		out549 => sig_1026,
		out550 => sig_1025,
		out552 => sig_1024,
		out558 => sig_1023,
		out559 => sig_1022,
		out563 => sig_1021,
		out566 => sig_1020,
		out572 => sig_1019,
		out573 => sig_1018,
		out576 => sig_1017,
		out577 => sig_1016,
		out581 => sig_1015,
		out582 => sig_1014,
		out590 => sig_1013,
		out591 => sig_1012,
		out592 => sig_1011,
		out593 => sig_1010,
		out595 => sig_1009,
		out611 => sig_1008,
		out619 => sig_1007,
		out638 => sig_1006,
		out643 => sig_1005,
		out644 => sig_1004,
		out645 => sig_1003,
		out646 => sig_1002,
		out648 => sig_1001,
		out650 => sig_1000,
		out652 => sig_999,
		out657 => sig_998,
		out659 => sig_997,
		out662 => sig_996,
		out677 => sig_995,
		out678 => sig_994,
		out679 => sig_993,
		out680 => sig_992,
		out682 => sig_991,
		out686 => sig_990,
		out692 => sig_989,
		out1218 => sig_988,
		out1219 => sig_987,
		out1220 => sig_986,
		out1221 => sig_985,
		out695 => sig_984,
		out697 => sig_983,
		out706 => sig_982,
		out719 => sig_981,
		out729 => sig_980,
		out744 => sig_979,
		out746 => sig_978,
		out748 => sig_977,
		out833 => sig_976,
		out834 => sig_975,
		out836 => sig_974,
		out837 => sig_973,
		out839 => sig_972,
		out840 => sig_971,
		out841 => sig_970,
		out844 => sig_969,
		out845 => sig_968,
		out846 => sig_967,
		out848 => sig_966,
		out850 => sig_965,
		out852 => sig_964,
		out854 => sig_963,
		out856 => sig_962,
		out858 => sig_961,
		out860 => sig_960,
		out863 => sig_959,
		out865 => sig_958,
		out866 => sig_957,
		out873 => sig_956,
		out877 => sig_955,
		out888 => sig_954,
		out891 => sig_953,
		out893 => sig_952,
		out895 => sig_951,
		out898 => sig_950,
		out900 => sig_949,
		out902 => sig_948,
		out903 => sig_947,
		out904 => sig_946,
		out905 => sig_945,
		out906 => sig_944,
		out907 => sig_943,
		out908 => sig_942,
		out909 => sig_941,
		out910 => sig_940,
		out912 => sig_939,
		out913 => sig_938,
		out914 => sig_937,
		out915 => sig_936,
		out917 => sig_935,
		out920 => sig_934,
		out921 => sig_933,
		out924 => sig_932,
		out934 => sig_931,
		out935 => sig_930,
		out937 => sig_929,
		out938 => sig_928,
		out940 => sig_927,
		out943 => sig_926,
		out945 => sig_925,
		out957 => sig_924,
		out958 => sig_923,
		out962 => sig_922,
		out968 => sig_921,
		out972 => sig_920,
		out973 => sig_919,
		out974 => sig_918,
		out975 => sig_917,
		out976 => sig_916,
		out980 => sig_915,
		out986 => sig_914,
		out988 => sig_913,
		out989 => sig_912,
		out990 => sig_911,
		out1004 => sig_910,
		out1008 => sig_909,
		out999 => sig_908,
		out1000 => sig_907,
		out1002 => sig_906,
		out1003 => sig_905,
		out1050 => sig_904,
		out1052 => sig_903,
		out1053 => sig_902,
		out1055 => sig_901,
		out1056 => sig_900,
		out1057 => sig_899,
		out1059 => sig_898,
		out1015 => sig_897,
		out1025 => sig_896,
		out1026 => sig_895,
		out1038 => sig_894,
		out1039 => sig_893,
		out1042 => sig_892,
		out1043 => sig_891,
		out1046 => sig_890,
		out1048 => sig_889,
		out1061 => sig_888,
		out1063 => sig_887,
		out1064 => sig_886,
		out1067 => sig_885,
		out1068 => sig_884,
		out1069 => sig_883,
		out1071 => sig_882,
		out1073 => sig_881,
		out1076 => sig_880,
		out1077 => sig_879,
		out1078 => sig_878,
		out1080 => sig_877,
		out1081 => sig_876,
		out1083 => sig_875,
		out1085 => sig_874,
		out1087 => sig_873,
		out1089 => sig_872,
		out1092 => sig_871,
		out1096 => sig_870,
		out1100 => sig_869,
		out1103 => sig_868,
		out1115 => sig_867,
		out1122 => sig_866,
		out1123 => sig_865,
		out1127 => sig_864,
		out1130 => sig_863,
		out1133 => sig_862,
		out1138 => sig_861,
		out1139 => sig_860,
		out1140 => sig_859,
		out1141 => sig_858,
		out1142 => sig_857,
		out1143 => sig_856,
		out1144 => sig_855,
		out1145 => sig_854,
		out1146 => sig_853,
		out1147 => sig_852,
		out1148 => sig_851,
		out1149 => sig_850,
		out1150 => sig_849,
		out1151 => sig_848,
		out1152 => sig_847,
		out1153 => sig_846,
		out1154 => sig_845,
		out1155 => sig_844,
		out1156 => sig_843,
		out1157 => sig_842,
		out1158 => sig_841,
		out1159 => sig_840,
		out1160 => sig_839,
		out1161 => sig_838,
		out1162 => sig_837,
		out1163 => sig_836,
		out1164 => sig_835,
		out1165 => sig_834,
		out1166 => sig_833,
		out1167 => sig_832,
		out1168 => sig_831,
		out1169 => sig_830,
		out1170 => sig_829,
		out1171 => sig_828,
		out1172 => sig_827,
		out1173 => sig_826,
		out1174 => sig_825,
		out1175 => sig_824,
		out1176 => sig_823,
		out1177 => sig_822,
		out1178 => sig_821,
		out1179 => sig_820,
		out1180 => sig_819,
		out1181 => sig_818,
		out1182 => sig_817,
		out1183 => sig_816,
		out1184 => sig_815,
		out1185 => sig_814,
		out1186 => sig_813,
		out1187 => sig_812,
		out1188 => sig_811,
		out1189 => sig_810,
		out1190 => sig_809,
		out1191 => sig_808,
		out1192 => sig_807,
		out1193 => sig_806,
		out1194 => sig_805,
		out1195 => sig_804,
		out1196 => sig_803,
		out1197 => sig_802,
		out1198 => sig_801,
		out1199 => sig_800,
		out1200 => sig_799,
		out1201 => sig_798,
		out1202 => sig_797,
		out1203 => sig_796,
		out1204 => sig_795,
		out1205 => sig_794,
		out1206 => sig_793,
		out1207 => sig_792,
		out1208 => sig_791,
		out1209 => sig_790,
		out1210 => sig_789,
		out1211 => sig_788,
		out1212 => sig_787,
		out1213 => sig_786,
		out1214 => sig_785,
		out1215 => sig_784,
		out1216 => sig_783,
		out1217 => sig_782
	);

	-- Behaviour of component 'and_757' model 'and'
	and_757 <=
		uppol1_apl1_53 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'or_758' model 'or'
	or_758 <=
		and_760 or
		and_759;

	-- Behaviour of component 'and_760' model 'and'
	and_760 <=
		uppol2_apl2_43 and
		sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305;

	-- Behaviour of component 'or_761' model 'or'
	or_761 <=
		sig_1304(31) & "0000000" or
		not_762 & "0000000";

	-- Behaviour of component 'not_762' model 'not'
	not_762 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'not_764' model 'not'
	not_764 <= not (
		logsch_nbh_57(31)
	);

	-- Behaviour of component 'not_766' model 'not'
	not_766 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'or_767' model 'or'
	or_767 <=
		sig_1303(31) & "0000000" or
		not_768 & "0000000";

	-- Behaviour of component 'mux_490' model 'mux'
	mux_490 <=
		(repeat(31, sig_895) and dec_rlt1);

	-- Behaviour of component 'and_744' model 'and'
	and_744 <=
		uppol1_apl1_53 and
		sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282;

	-- Behaviour of component 'not_746' model 'not'
	not_746 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'or_747' model 'or'
	or_747 <=
		and_749 or
		and_748;

	-- Behaviour of component 'and_748' model 'and'
	and_748 <=
		"00000000000000000011000000000000" and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'not_751' model 'not'
	not_751 <= not (
		logsch_nbh_57(31)
	);

	-- Behaviour of component 'or_752' model 'or'
	or_752 <=
		and_754 or
		and_753;

	-- Behaviour of component 'and_753' model 'and'
	and_753 <=
		sig_1307(31 downto 0) and
		sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301;

	-- Behaviour of component 'or_755' model 'or'
	or_755 <=
		and_757 or
		and_756;

	-- Behaviour of component 'or_714' model 'or'
	or_714 <=
		and_716 or
		and_715;

	-- Behaviour of component 'and_715' model 'and'
	and_715 <=
		"11111111111111111101000000000000" and
		sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301;

	-- Behaviour of component 'and_723' model 'and'
	and_723 <=
		sig_1302(31 downto 0) and
		sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31);

	-- Behaviour of component 'and_727' model 'and'
	and_727 <=
		sig_1290(25 downto 0) & uppol1_wd2_51(5 downto 0) and
		not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728 & not_728;

	-- Behaviour of component 'not_728' model 'not'
	not_728 <= not (
		sig_1281(31)
	);

	-- Behaviour of component 'and_735' model 'and'
	and_735 <=
		uppol1_wd3_52 and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'or_742' model 'or'
	or_742 <=
		and_744 or
		and_743;

	-- Behaviour of component 'and_743' model 'and'
	and_743 <=
		sig_1307(31 downto 0) and
		sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301;

	-- Behaviour of component 'mux_484' model 'mux'
	mux_484 <=
		(repeat(32, sig_993) and uppol1_apl1_53);

	-- Behaviour of component 'mux_486' model 'mux'
	mux_486 <=
		(repeat(32, sig_1015) and uppol2_apl2_43);

	-- Behaviour of component 'mux_488' model 'mux'
	mux_488 <=
		(repeat(31, sig_1133) and dec_rlt);

	-- Behaviour of component 'mux_480' model 'mux'
	mux_480 <=
		(repeat(32, sig_1015) and logsch_nbh_57);

	-- Behaviour of component 'mux_476' model 'mux'
	mux_476 <=
		(repeat(32, sig_1033) and logscl_nbl_27);

	-- Behaviour of component 'mux_472' model 'mux'
	mux_472 <=
		(repeat(31, sig_954) and rh(30 downto 0));

	-- Behaviour of component 'mux_474' model 'mux'
	mux_474 <=
		(repeat(31, sig_1257) and dec_rh1);

	-- Behaviour of component 'mux_470' model 'mux'
	mux_470 <=
		(repeat(32, sig_1027) and uppol2_apl2_43);

	-- Behaviour of component 'mux_468' model 'mux'
	mux_468 <=
		(repeat(32, sig_1059) and uppol1_apl1_53);

	-- Behaviour of component 'mux_460' model 'mux'
	mux_460 <=
		(repeat(32, sig_954) and dec_ph);

	-- Behaviour of component 'mux_462' model 'mux'
	mux_462 <=
		(repeat(32, sig_1257) and dec_ph1);

	-- Behaviour of component 'mux_456' model 'mux'
	mux_456 <=
		(repeat(64, sig_1133) and sig_1298) or
		(repeat(64, sig_1154) and sig_1303) or
		(repeat(64, sig_1241) and sig_1290) or
		(repeat(64, sig_868) and sig_1281) or
		(repeat(64, sig_895) and sig_1287) or
		(repeat(64, sig_926) and sig_1289);

	-- Behaviour of component 'mux_458' model 'mux'
	mux_458 <=
		(repeat(32, sig_966) and or_710) or
		(repeat(32, sig_976) and or_705);

	-- Behaviour of component 'mux_448' model 'mux'
	mux_448 <=
		(repeat(32, sig_901) and sig_1298(31 downto 0));

	-- Behaviour of component 'mux_434' model 'mux'
	mux_434 <=
		(repeat(32, sig_997) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_697) or
		(repeat(32, sig_1153) and sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & or_636) or
		(repeat(32, sig_1257) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_627) or
		(repeat(32, sig_895) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_740);

	-- Behaviour of component 'mux_438' model 'mux'
	mux_438 <=
		(repeat(32, sig_911) and sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31 downto 7)) or
		(repeat(32, sig_1061) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 7));

	-- Behaviour of component 'mux_440' model 'mux'
	mux_440 <=
		(repeat(32, sig_1038) and and_681) or
		(repeat(32, sig_1099) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1107) and or_648) or
		(repeat(32, sig_935) and and_724) or
		(repeat(32, sig_1034) and or_685);

	-- Behaviour of component 'mux_430' model 'mux'
	mux_430 <=
		(repeat(32, sig_1149) and sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31 downto 8)) or
		(repeat(32, sig_1256) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31 downto 8));

	-- Behaviour of component 'mux_432' model 'mux'
	mux_432 <=
		(repeat(32, sig_927) and sig_1288(31 downto 0)) or
		(repeat(32, sig_908) and or_737) or
		(repeat(32, sig_1133) and sig_1286) or
		(repeat(32, sig_955) and or_717) or
		(repeat(32, sig_1142) and or_641) or
		(repeat(32, sig_1166) and or_631) or
		(repeat(32, sig_961) and or_714) or
		(repeat(32, sig_1022) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1091) and or_657) or
		(repeat(32, sig_904) and or_747) or
		(repeat(32, sig_879) and or_758);

	-- Behaviour of component 'mux_424' model 'mux'
	mux_424 <=
		(repeat(32, sig_1072) and or_666) or
		(repeat(32, sig_1133) and sig_1289(31 downto 0)) or
		(repeat(32, sig_1142) and or_638) or
		(repeat(32, sig_869) and sig_1298(31 downto 0)) or
		(repeat(32, sig_874) and and_763) or
		(repeat(32, sig_904) and and_750);

	-- Behaviour of component 'mux_426' model 'mux'
	mux_426 <=
		(repeat(32, sig_916) and or_734) or
		(repeat(32, sig_893) and or_742) or
		(repeat(32, sig_1093) and or_654) or
		(repeat(32, sig_927) and or_726) or
		(repeat(32, sig_1101) and or_651) or
		(repeat(32, sig_1133) and or_644) or
		(repeat(32, sig_954) and or_720) or
		(repeat(32, sig_1023) and or_688) or
		(repeat(32, sig_1082) and or_663) or
		(repeat(32, sig_885) and or_752) or
		(repeat(32, sig_882) and or_755) or
		(repeat(32, sig_865) and or_769);

	-- Behaviour of component 'mux_422' model 'mux'
	mux_422 <=
		(repeat(32, sig_895) and sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31 downto 7)) or
		(repeat(32, sig_1153) and sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31 downto 7));

	-- Behaviour of component 'mux_416' model 'mux'
	mux_416 <=
		(repeat(64, sig_868) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 0)) or
		(repeat(64, sig_1260) and sig_1298) or
		(repeat(64, sig_1198) and sig_1289);

	-- Behaviour of component 'mux_414' model 'mux'
	mux_414 <=
		(repeat(64, sig_868) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31 downto 0)) or
		(repeat(64, sig_1260) and sig_1289) or
		(repeat(64, sig_1198) and sig_1298);

	-- Behaviour of component 'mux_406' model 'mux'
	mux_406 <=
		(repeat(64, sig_955) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31 downto 0)) or
		(repeat(64, sig_1066) and sig_1289) or
		(repeat(64, sig_1145) and sig_1298);

	-- Behaviour of component 'mux_400' model 'mux'
	mux_400 <=
		(repeat(32, sig_1252) and "00000000000000000000000000001100") or
		(repeat(32, sig_1172) and "00000000000000000000000000000000") or
		(repeat(32, sig_1278) and "00000000000000000000000011111111") or
		(repeat(32, sig_1254) and "00000000000000000011110010010000") or
		(repeat(32, sig_1243) and "00000000000000000000000011010100") or
		(repeat(32, sig_1196) and "00000000000000000000010110101000") or
		(repeat(32, sig_1257) and dec_ph2) or
		(repeat(32, sig_1262) and dec_del_dltx_reg1) or
		(repeat(32, sig_1273) and delay_dhx_reg0) or
		(repeat(32, sig_1163) and "00000000000000000000000000000000") or
		(repeat(32, sig_1159) and quantl_detl_17) or
		(repeat(32, sig_1147) and "11111111111111111111110110010000") or
		(repeat(32, sig_1142) and "00000000000000000000000000000000") or
		(repeat(32, sig_1133) and dec_ah2) or
		(repeat(32, sig_1119) and "11111111111111111111001101101100") or
		(repeat(32, sig_1101) and "00000000000000000000000000000000") or
		(repeat(32, sig_1099) and sig_1316) or
		(repeat(32, sig_1065) and "00000000000000000000111011011100") or
		(repeat(32, sig_1062) and "00000000000000000000000001111111") or
		(repeat(32, sig_1049) and "11111111111111111111110010111000") or
		(repeat(32, sig_1042) and "00000000000000000000000000000000") or
		(repeat(32, sig_1040) and "00000000000000000000000000000000") or
		(repeat(32, sig_1038) and "00000000000000000000000000000000") or
		(repeat(32, sig_1034) and "00000000000000000000000000000000") or
		(repeat(32, sig_1033) and "00000000000000000000000000000000") or
		(repeat(32, sig_1009) and "11111111111111111111111111010100") or
		(repeat(32, sig_1003) and "00000000000000000000000000000000") or
		(repeat(32, sig_997) and ph2) or
		(repeat(32, sig_970) and "00000000000000000000000000110000") or
		(repeat(32, sig_930) and "00000000000000000000000010000000") or
		(repeat(32, sig_928) and delay_dhx_reg1) or
		(repeat(32, sig_923) and delay_dltx_reg1) or
		(repeat(32, sig_922) and delay_dltx_reg0) or
		(repeat(32, sig_912) and dec_del_dltx_reg0) or
		(repeat(32, sig_909) and sig_1309) or
		(repeat(32, sig_889) and "00000000000000000000000000000000") or
		(repeat(32, sig_883) and "00000000000000000000000000000000") or
		(repeat(32, sig_879) and "00000000000000000000000000000000") or
		(repeat(32, sig_1200) and dec_del_dhx_reg0);

	-- Behaviour of component 'mux_402' model 'mux'
	mux_402 <=
		(repeat(64, sig_1031) and "0000000000000000000000000000000000000000000000000000000000001000") or
		(repeat(64, sig_1015) and logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16 downto 11)) or
		(repeat(64, sig_1108) and logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27) or
		(repeat(64, sig_1045) and ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih(31) & ih) or
		(repeat(64, sig_1143) and logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57) or
		(repeat(64, sig_1168) and uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43) or
		(repeat(64, sig_1069) and "0000000000000000000000000000000000000000000000000000000000001010") or
		(repeat(64, sig_1102) and uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53) or
		(repeat(64, sig_954) and rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl);

	-- Behaviour of component 'mux_403' model 'mux'
	mux_403 <=
		(repeat(64, sig_954) and rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh) or
		(repeat(64, sig_1108) and "0000000000000000000000000000000000000000000000000100100000000000") or
		(repeat(64, sig_962) and "1111111111111111111111111111111111111111111111111101000000000000") or
		(repeat(64, sig_1143) and "0000000000000000000000000000000000000000000000000101100000000000") or
		(repeat(64, sig_1167) and "0000000000000000000000000000000000000000000000000011000000000000") or
		(repeat(64, sig_1044) and "0000000000000000000000000000000000000000000000000000000000000001") or
		(repeat(64, sig_1068) and sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5) & sig_1302(5 downto 0)) or
		(repeat(64, sig_1103) and uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52);

	-- Behaviour of component 'mux_404' model 'mux'
	mux_404 <=
		(repeat(64, sig_955) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 0)) or
		(repeat(64, sig_1066) and sig_1298) or
		(repeat(64, sig_1145) and sig_1289);

	-- Behaviour of component 'mux_395' model 'mux'
	mux_395 <=
		(repeat(64, sig_1031) and logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16) & logscl_nbl_27(16 downto 11)) or
		(repeat(64, sig_1029) and "0000000000000000000000000000000000000000000000000011110000000000") or
		(repeat(64, sig_1135) and uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51) or
		(repeat(64, sig_1045) and abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3) or
		(repeat(64, sig_1143) and logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57(31) & logsch_nbh_57) or
		(repeat(64, sig_1168) and uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43) or
		(repeat(64, sig_1069) and logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16) & logsch_nbh_57(16 downto 11)) or
		(repeat(64, sig_1103) and uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53) or
		(repeat(64, sig_1108) and logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27(31) & logscl_nbl_27) or
		(repeat(64, sig_964) and xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh(31) & xh) or
		(repeat(64, sig_959) and xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl(31) & xl) or
		(repeat(64, sig_957) and encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46 downto 0)) or
		(repeat(64, sig_951) and augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132) or
		(repeat(64, sig_898) and quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19) or
		(repeat(64, sig_881) and quantl_wd_20);

	-- Behaviour of component 'mux_396' model 'mux'
	mux_396 <=
		(repeat(64, sig_1045) and encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69) or
		(repeat(64, sig_1029) and uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43) or
		(repeat(64, sig_1135) and "0000000000000000000000000000000000000000000000000000000011000000") or
		(repeat(64, sig_1068) and "0000000000000000000000000000000000000000000000000000000000000001") or
		(repeat(64, sig_1143) and "0000000000000000000000000000000000000000000000000101100000000000") or
		(repeat(64, sig_1167) and "0000000000000000000000000000000000000000000000000011000000000000") or
		(repeat(64, sig_1094) and sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31 downto 0)) or
		(repeat(64, sig_1102) and uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52(31) & uppol1_wd3_52) or
		(repeat(64, sig_1108) and "0000000000000000000000000000000000000000000000000100100000000000") or
		(repeat(64, sig_976) and eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh) or
		(repeat(64, sig_966) and el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el) or
		(repeat(64, sig_964) and sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh) or
		(repeat(64, sig_962) and "1111111111111111111111111111111111111111111111111101000000000000") or
		(repeat(64, sig_959) and sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl) or
		(repeat(64, sig_957) and encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46 downto 0)) or
		(repeat(64, sig_951) and "0000000000000000000000000000000000000000000000000000000001100011") or
		(repeat(64, sig_898) and "0000000000000000000000000000000000000000000000000000000000011101") or
		(repeat(64, sig_881) and "00000000000000000000000000000000" & quantl_decis_21);

	-- Behaviour of component 'mux_397' model 'mux'
	mux_397 <=
		(repeat(64, sig_1257) and dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1(31) & dec_ah1) or
		(repeat(64, sig_1253) and tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10(31) & tqmf_reg10) or
		(repeat(64, sig_1275) and dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh) or
		(repeat(64, sig_1261) and tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21(31) & tqmf_reg21) or
		(repeat(64, sig_1241) and tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2(31) & tqmf_reg2) or
		(repeat(64, sig_1195) and tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6(31) & tqmf_reg6) or
		(repeat(64, sig_1262) and dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1(31) & dec_del_bpl_reg1) or
		(repeat(64, sig_1265) and dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt) or
		(repeat(64, sig_1270) and delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0) or
		(repeat(64, sig_1175) and tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22(31) & tqmf_reg22) or
		(repeat(64, sig_1174) and dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5) or
		(repeat(64, sig_1160) and dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4) or
		(repeat(64, sig_1153) and rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1(30) & rh1 & '0') or
		(repeat(64, sig_1146) and accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8(31) & accumd_reg8) or
		(repeat(64, sig_1136) and dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt(31) & dec_plt) or
		(repeat(64, sig_1125) and delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5) or
		(repeat(64, sig_1118) and accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6(31) & accumd_reg6) or
		(repeat(64, sig_1115) and delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5) or
		(repeat(64, sig_1085) and dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt) or
		(repeat(64, sig_1064) and accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5(31) & accumc_reg5) or
		(repeat(64, sig_1059) and accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4(31) & accumd_reg4) or
		(repeat(64, sig_1053) and dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4) or
		(repeat(64, sig_1048) and tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14(31) & tqmf_reg14) or
		(repeat(64, sig_1042) and delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2(31) & delay_bpl_reg2) or
		(repeat(64, sig_1040) and delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3(31) & delay_bpl_reg3) or
		(repeat(64, sig_1035) and tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17(31) & tqmf_reg17) or
		(repeat(64, sig_1027) and accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1(31) & accumc_reg1) or
		(repeat(64, sig_1023) and ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph) or
		(repeat(64, sig_1016) and tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9(31) & tqmf_reg9) or
		(repeat(64, sig_1008) and accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10(31) & accumd_reg10) or
		(repeat(64, sig_997) and ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1(31) & ah1) or
		(repeat(64, sig_973) and dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh) or
		(repeat(64, sig_969) and tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18(31) & tqmf_reg18) or
		(repeat(64, sig_961) and accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0(31) & accumd_reg0) or
		(repeat(64, sig_955) and xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd(31) & xd) or
		(repeat(64, sig_954) and dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph) or
		(repeat(64, sig_931) and accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7(31) & accumc_reg7) or
		(repeat(64, sig_927) and rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2(30) & rh2 & '0') or
		(repeat(64, sig_923) and delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1(31) & delay_bpl_reg1) or
		(repeat(64, sig_922) and delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0) or
		(repeat(64, sig_921) and tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13(31) & tqmf_reg13) or
		(repeat(64, sig_914) and dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2(30) & dec_rlt2 & '0') or
		(repeat(64, sig_911) and dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1(30) & dec_rlt1 & '0') or
		(repeat(64, sig_887) and accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9(31) & accumc_reg9) or
		(repeat(64, sig_885) and accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3(31) & accumc_reg3) or
		(repeat(64, sig_872) and dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0) or
		(repeat(64, sig_868) and tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1(31) & tqmf_reg1) or
		(repeat(64, sig_866) and tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5(31) & tqmf_reg5) or
		(repeat(64, sig_865) and accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2(31) & accumd_reg2) or
		(repeat(64, sig_864) and delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1) or
		(repeat(64, sig_861) and dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2) or
		(repeat(64, sig_1200) and dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0);

	-- Behaviour of component 'mux_398' model 'mux'
	mux_398 <=
		(repeat(32, sig_1147) and "00000000000000000000000000110000") or
		(repeat(32, sig_1133) and dec_plt1) or
		(repeat(32, sig_1153) and ah1) or
		(repeat(32, sig_1242) and "11111111111111111111111111010100") or
		(repeat(32, sig_1196) and "00000000000000000000000010000000") or
		(repeat(32, sig_1254) and "00000000000000000000111011011100") or
		(repeat(32, sig_1268) and "00000000000000000000000000000000") or
		(repeat(32, sig_1271) and "00000000000000000000000011111111") or
		(repeat(32, sig_1119) and "11111111111111111111110010111000") or
		(repeat(32, sig_1086) and "00000000000000000000000000000000") or
		(repeat(32, sig_1065) and "00000000000000000011110010010000") or
		(repeat(32, sig_1049) and "11111111111111111111001101101100") or
		(repeat(32, sig_1036) and "00000000000000000000000000000000") or
		(repeat(32, sig_1023) and ph1) or
		(repeat(32, sig_1017) and "00000000000000000000000000000000") or
		(repeat(32, sig_1007) and "00000000000000000000000000001100") or
		(repeat(32, sig_1000) and "00000000000000000000000000000000") or
		(repeat(32, sig_974) and "00000000000000000000000000000000") or
		(repeat(32, sig_970) and "11111111111111111111110110010000") or
		(repeat(32, sig_960) and "00000000000000000000000011010100") or
		(repeat(32, sig_954) and dec_ph1) or
		(repeat(32, sig_930) and "00000000000000000000010110101000") or
		(repeat(32, sig_927) and ah2) or
		(repeat(32, sig_914) and dec_al2) or
		(repeat(32, sig_911) and dec_al1) or
		(repeat(32, sig_895) and dec_plt2) or
		(repeat(32, sig_890) and "00000000000000000000000000000000") or
		(repeat(32, sig_871) and "00000000000000000000000000000000") or
		(repeat(32, sig_863) and "00000000000000000000000000000000") or
		(repeat(32, sig_862) and dec_del_dhx_reg1);

	-- Behaviour of component 'mux_399' model 'mux'
	mux_399 <=
		(repeat(64, sig_1257) and dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph(31) & dec_ph) or
		(repeat(64, sig_1253) and tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11(31) & tqmf_reg11) or
		(repeat(64, sig_1277) and delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2(31) & delay_bph_reg2) or
		(repeat(64, sig_1261) and tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20(31) & tqmf_reg20) or
		(repeat(64, sig_1241) and tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3(31) & tqmf_reg3) or
		(repeat(64, sig_1195) and tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7(31) & tqmf_reg7) or
		(repeat(64, sig_1263) and dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt) or
		(repeat(64, sig_1266) and dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3(31) & dec_del_bpl_reg3) or
		(repeat(64, sig_1272) and dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh) or
		(repeat(64, sig_1175) and tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23(31) & tqmf_reg23) or
		(repeat(64, sig_1162) and dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh) or
		(repeat(64, sig_1159) and sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312(31) & sig_1312) or
		(repeat(64, sig_1155) and delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0(31) & delay_bph_reg0) or
		(repeat(64, sig_1146) and accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8(31) & accumc_reg8) or
		(repeat(64, sig_1140) and dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3(31) & dec_del_bph_reg3) or
		(repeat(64, sig_1133) and dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2(30) & dec_rh2 & '0') or
		(repeat(64, sig_1125) and delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0(31) & delay_bpl_reg0) or
		(repeat(64, sig_1122) and dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5(31) & dec_del_bpl_reg5) or
		(repeat(64, sig_1118) and accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6(31) & accumc_reg6) or
		(repeat(64, sig_1104) and dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5(31) & dec_del_bph_reg5) or
		(repeat(64, sig_1100) and detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl(31) & detl) or
		(repeat(64, sig_1086) and delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5(31) & delay_bpl_reg5) or
		(repeat(64, sig_1064) and accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5(31) & accumd_reg5) or
		(repeat(64, sig_1061) and nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl(31) & nbl) or
		(repeat(64, sig_1059) and accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4(31) & accumc_reg4) or
		(repeat(64, sig_1054) and dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0(31) & dec_del_bpl_reg0) or
		(repeat(64, sig_1048) and tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15(31) & tqmf_reg15) or
		(repeat(64, sig_1041) and dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt) or
		(repeat(64, sig_1037) and dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2(31) & dec_del_bpl_reg2) or
		(repeat(64, sig_1036) and delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4(31) & delay_bpl_reg4) or
		(repeat(64, sig_1035) and tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16(31) & tqmf_reg16) or
		(repeat(64, sig_1032) and dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4(31) & dec_del_bpl_reg4) or
		(repeat(64, sig_1027) and accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1(31) & accumd_reg1) or
		(repeat(64, sig_1023) and ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2(31) & ah2) or
		(repeat(64, sig_1016) and tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8(31) & tqmf_reg8) or
		(repeat(64, sig_1015) and dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4(31) & dec_del_bph_reg4) or
		(repeat(64, sig_1008) and accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10(31) & accumc_reg10) or
		(repeat(64, sig_1002) and delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4(31) & delay_bph_reg4) or
		(repeat(64, sig_997) and ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph(31) & ph) or
		(repeat(64, sig_969) and tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19(31) & tqmf_reg19) or
		(repeat(64, sig_961) and accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0(31) & accumc_reg0) or
		(repeat(64, sig_955) and xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs(31) & xs) or
		(repeat(64, sig_954) and dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2(31) & dec_ah2) or
		(repeat(64, sig_932) and dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0(31) & dec_del_bph_reg0) or
		(repeat(64, sig_931) and accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7(31) & accumd_reg7) or
		(repeat(64, sig_927) and delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1(31) & delay_bph_reg1) or
		(repeat(64, sig_921) and tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12(31) & tqmf_reg12) or
		(repeat(64, sig_914) and dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl(31) & dec_detl) or
		(repeat(64, sig_895) and dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth(31) & dec_deth) or
		(repeat(64, sig_904) and dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2(31) & dec_del_bph_reg2) or
		(repeat(64, sig_887) and accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9(31) & accumd_reg9) or
		(repeat(64, sig_885) and accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3(31) & accumd_reg3) or
		(repeat(64, sig_882) and delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5(31) & delay_bph_reg5) or
		(repeat(64, sig_880) and delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3(31) & delay_bph_reg3) or
		(repeat(64, sig_869) and deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth(31) & deth) or
		(repeat(64, sig_868) and tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0(31) & tqmf_reg0) or
		(repeat(64, sig_866) and tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4(31) & tqmf_reg4) or
		(repeat(64, sig_865) and accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2(31) & accumc_reg2) or
		(repeat(64, sig_862) and dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1(31) & dec_del_bph_reg1);

	-- Behaviour of component 'mux_383' model 'mux'
	mux_383 <=
		(repeat(6, sig_1015) and sig_1285(5 downto 0)) or
		(repeat(6, sig_1068) and sig_1307(5 downto 0));

	-- Behaviour of component 'mux_385' model 'mux'
	mux_385 <=
		(repeat(7, sig_1139) and "1100011") or
		(repeat(7, sig_1047) and "0000110") or
		(repeat(7, sig_1182) and "0000101") or
		(repeat(7, sig_1183) and "0001000") or
		(repeat(7, sig_1214) and "0001010") or
		(repeat(7, sig_1192) and "0000010") or
		(repeat(7, sig_1189) and "0000011") or
		(repeat(7, sig_1187) and "0000111") or
		(repeat(7, sig_1025) and "0001001") or
		(repeat(7, sig_1019) and "0000001") or
		(repeat(7, sig_999) and "0000100") or
		(repeat(7, sig_860) and "1100010") or
		(repeat(7, sig_859) and "1100001") or
		(repeat(7, sig_858) and "1100000") or
		(repeat(7, sig_857) and "1011111") or
		(repeat(7, sig_856) and "1011110") or
		(repeat(7, sig_855) and "1011101") or
		(repeat(7, sig_854) and "1011100") or
		(repeat(7, sig_853) and "1011011") or
		(repeat(7, sig_852) and "1011010") or
		(repeat(7, sig_851) and "1011001") or
		(repeat(7, sig_850) and "1011000") or
		(repeat(7, sig_849) and "1010111") or
		(repeat(7, sig_848) and "1010110") or
		(repeat(7, sig_847) and "1010101") or
		(repeat(7, sig_846) and "1010100") or
		(repeat(7, sig_845) and "1010011") or
		(repeat(7, sig_844) and "1010010") or
		(repeat(7, sig_843) and "1010001") or
		(repeat(7, sig_842) and "1010000") or
		(repeat(7, sig_841) and "1001111") or
		(repeat(7, sig_840) and "1001110") or
		(repeat(7, sig_839) and "1001101") or
		(repeat(7, sig_838) and "1001100") or
		(repeat(7, sig_837) and "1001011") or
		(repeat(7, sig_836) and "1001010") or
		(repeat(7, sig_835) and "1001001") or
		(repeat(7, sig_834) and "1001000") or
		(repeat(7, sig_833) and "1000111") or
		(repeat(7, sig_832) and "1000110") or
		(repeat(7, sig_831) and "1000101") or
		(repeat(7, sig_830) and "1000100") or
		(repeat(7, sig_829) and "1000011") or
		(repeat(7, sig_828) and "1000010") or
		(repeat(7, sig_827) and "1000001") or
		(repeat(7, sig_826) and "1000000") or
		(repeat(7, sig_825) and "0111111") or
		(repeat(7, sig_824) and "0111110") or
		(repeat(7, sig_823) and "0111101") or
		(repeat(7, sig_822) and "0111100") or
		(repeat(7, sig_821) and "0111011") or
		(repeat(7, sig_820) and "0111010") or
		(repeat(7, sig_819) and "0111001") or
		(repeat(7, sig_818) and "0111000") or
		(repeat(7, sig_817) and "0110111") or
		(repeat(7, sig_816) and "0110110") or
		(repeat(7, sig_815) and "0110101") or
		(repeat(7, sig_814) and "0110100") or
		(repeat(7, sig_813) and "0110011") or
		(repeat(7, sig_812) and "0110010") or
		(repeat(7, sig_811) and "0110001") or
		(repeat(7, sig_810) and "0110000") or
		(repeat(7, sig_809) and "0101111") or
		(repeat(7, sig_808) and "0101110") or
		(repeat(7, sig_807) and "0101101") or
		(repeat(7, sig_806) and "0101100") or
		(repeat(7, sig_805) and "0101011") or
		(repeat(7, sig_804) and "0101010") or
		(repeat(7, sig_803) and "0101001") or
		(repeat(7, sig_802) and "0101000") or
		(repeat(7, sig_801) and "0100111") or
		(repeat(7, sig_800) and "0100110") or
		(repeat(7, sig_799) and "0100101") or
		(repeat(7, sig_798) and "0100100") or
		(repeat(7, sig_797) and "0100011") or
		(repeat(7, sig_796) and "0100010") or
		(repeat(7, sig_795) and "0100001") or
		(repeat(7, sig_794) and "0100000") or
		(repeat(7, sig_793) and "0011111") or
		(repeat(7, sig_792) and "0011110") or
		(repeat(7, sig_791) and "0011101") or
		(repeat(7, sig_790) and "0011100") or
		(repeat(7, sig_789) and "0011011") or
		(repeat(7, sig_788) and "0011010") or
		(repeat(7, sig_787) and "0011001") or
		(repeat(7, sig_786) and "0011000") or
		(repeat(7, sig_785) and "0010111") or
		(repeat(7, sig_784) and "0010110") or
		(repeat(7, sig_783) and "0010101") or
		(repeat(7, sig_782) and "0010100") or
		(repeat(7, sig_988) and "0010011") or
		(repeat(7, sig_987) and "0010010") or
		(repeat(7, sig_986) and "0010001") or
		(repeat(7, sig_985) and "0010000") or
		(repeat(7, sig_1205) and "0001111") or
		(repeat(7, sig_1204) and "0001110") or
		(repeat(7, sig_1203) and "0001101") or
		(repeat(7, sig_1202) and "0001100") or
		(repeat(7, sig_1201) and "0001011");

	-- Behaviour of component 'mux_390' model 'mux'
	mux_390 <=
		(repeat(64, sig_1133) and filtep_pl_14) or
		(repeat(64, sig_1099) and logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28(31) & logscl_wd_28) or
		(repeat(64, sig_1260) and encode_xa_67) or
		(repeat(64, sig_1145) and decode_xa1_100) or
		(repeat(64, sig_1231) and upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2(31) & upzero_wd2) or
		(repeat(64, sig_1198) and encode_xb_68) or
		(repeat(64, sig_1153) and sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl(31) & sl) or
		(repeat(64, sig_1169) and filtez_zl) or
		(repeat(64, sig_1257) and dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh(31) & dec_sh) or
		(repeat(64, sig_1097) and filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46 downto 15)) or
		(repeat(64, sig_1090) and augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6) & augh_main_i_132(6 downto 0)) or
		(repeat(64, sig_1084) and dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl(31) & dl) or
		(repeat(64, sig_1066) and decode_xa2_101) or
		(repeat(64, sig_1022) and uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42) or
		(repeat(64, sig_997) and sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh(31) & sh) or
		(repeat(64, sig_957) and encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46) & encode_xa_67(46 downto 0)) or
		(repeat(64, sig_950) and augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31 downto 1)) or
		(repeat(64, sig_935) and dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt) or
		(repeat(64, sig_895) and dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl) or
		(repeat(64, sig_893) and dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh) or
		(repeat(64, sig_901) and quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19(31) & quantl_mil_19) or
		(repeat(64, sig_874) and dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh) or
		(repeat(64, sig_869) and logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58);

	-- Behaviour of component 'mux_391' model 'mux'
	mux_391 <=
		(repeat(64, sig_1089) and "0000000000000000000000000000000000000000000000000000000000000001") or
		(repeat(64, sig_1084) and dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl(31) & dec_sl) or
		(repeat(64, sig_1257) and dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh(31) & dec_dh) or
		(repeat(64, sig_1096) and filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45 downto 14)) or
		(repeat(64, sig_1231) and upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3(31) & upzero_wd3) or
		(repeat(64, sig_1194) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 0)) or
		(repeat(64, sig_1099) and sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314(31) & sig_1314) or
		(repeat(64, sig_1133) and sig_1304) or
		(repeat(64, sig_1153) and dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt(31) & dlt) or
		(repeat(64, sig_1022) and sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38) & sig_1304(38 downto 7)) or
		(repeat(64, sig_997) and dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh(31) & dh) or
		(repeat(64, sig_957) and encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46) & encode_xb_68(46 downto 0)) or
		(repeat(64, sig_935) and szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl(31) & szl) or
		(repeat(64, sig_895) and dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt) or
		(repeat(64, sig_869) and sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308);

	-- Behaviour of component 'mux_376' model 'mux'
	mux_376 <=
		(repeat(7, sig_1222) and "1001111") or
		(repeat(7, sig_1220) and "1000001") or
		(repeat(7, sig_1211) and "0100110") or
		(repeat(7, sig_1223) and "1010000") or
		(repeat(7, sig_1212) and "1000110") or
		(repeat(7, sig_1210) and "0000111") or
		(repeat(7, sig_1224) and "0011111") or
		(repeat(7, sig_1217) and "0000100") or
		(repeat(7, sig_1216) and "0001100") or
		(repeat(7, sig_1219) and "0111000") or
		(repeat(7, sig_1218) and "1001001") or
		(repeat(7, sig_1230) and "1000000") or
		(repeat(7, sig_1229) and "0100001") or
		(repeat(7, sig_1228) and "1011000") or
		(repeat(7, sig_1245) and "1000111") or
		(repeat(7, sig_1244) and "1010111") or
		(repeat(7, sig_1247) and "0101001") or
		(repeat(7, sig_1246) and "0010101") or
		(repeat(7, sig_1250) and "0000011") or
		(repeat(7, sig_1249) and "0010110") or
		(repeat(7, sig_1248) and "0010111") or
		(repeat(7, sig_1251) and "0001110") or
		(repeat(7, sig_1236) and "0001011") or
		(repeat(7, sig_1235) and "1010001") or
		(repeat(7, sig_1239) and "0011000") or
		(repeat(7, sig_1238) and "1010010") or
		(repeat(7, sig_1237) and "1011010") or
		(repeat(7, sig_1208) and "1011011") or
		(repeat(7, sig_1207) and "1011001") or
		(repeat(7, sig_1206) and "0010010") or
		(repeat(7, sig_1234) and "1001000") or
		(repeat(7, sig_1233) and "1010100") or
		(repeat(7, sig_1180) and "1001011") or
		(repeat(7, sig_1179) and "0101011") or
		(repeat(7, sig_1178) and "1001101") or
		(repeat(7, sig_1177) and "1000101") or
		(repeat(7, sig_1185) and "1000100") or
		(repeat(7, sig_1184) and "0110101") or
		(repeat(7, sig_1181) and "0001000") or
		(repeat(7, sig_1188) and "0100100") or
		(repeat(7, sig_1186) and "0100000") or
		(repeat(7, sig_1190) and "0110000") or
		(repeat(7, sig_1191) and "0011001") or
		(repeat(7, sig_1193) and "0000110") or
		(repeat(7, sig_1157) and "0010001") or
		(repeat(7, sig_1156) and "0001111") or
		(repeat(7, sig_1137) and "1010101") or
		(repeat(7, sig_1123) and "1010110") or
		(repeat(7, sig_1120) and "0110011") or
		(repeat(7, sig_1117) and "0111110") or
		(repeat(7, sig_1109) and "0000101") or
		(repeat(7, sig_1080) and "1100011") or
		(repeat(7, sig_1079) and "1100010") or
		(repeat(7, sig_1078) and "1100001") or
		(repeat(7, sig_1077) and "1100000") or
		(repeat(7, sig_1076) and "1011111") or
		(repeat(7, sig_1075) and "1011110") or
		(repeat(7, sig_1074) and "1011101") or
		(repeat(7, sig_1073) and "1011100") or
		(repeat(7, sig_1055) and "0100111") or
		(repeat(7, sig_1046) and "0110010") or
		(repeat(7, sig_1039) and "0011101") or
		(repeat(7, sig_1018) and "1000010") or
		(repeat(7, sig_1013) and "0011110") or
		(repeat(7, sig_1012) and "0110111") or
		(repeat(7, sig_991) and "0000001") or
		(repeat(7, sig_972) and "0100011") or
		(repeat(7, sig_971) and "0011010") or
		(repeat(7, sig_968) and "0111100") or
		(repeat(7, sig_967) and "0110110") or
		(repeat(7, sig_952) and "0101000") or
		(repeat(7, sig_948) and "0111011") or
		(repeat(7, sig_947) and "1000011") or
		(repeat(7, sig_946) and "0111111") or
		(repeat(7, sig_945) and "0111001") or
		(repeat(7, sig_944) and "1001010") or
		(repeat(7, sig_943) and "1001100") or
		(repeat(7, sig_942) and "0101101") or
		(repeat(7, sig_941) and "1010011") or
		(repeat(7, sig_940) and "0101110") or
		(repeat(7, sig_939) and "0110100") or
		(repeat(7, sig_938) and "0100010") or
		(repeat(7, sig_937) and "0010100") or
		(repeat(7, sig_933) and "0101111") or
		(repeat(7, sig_929) and "0010011") or
		(repeat(7, sig_924) and "0101100") or
		(repeat(7, sig_919) and "0000010") or
		(repeat(7, sig_918) and "0011100") or
		(repeat(7, sig_917) and "0001010") or
		(repeat(7, sig_907) and "0010000") or
		(repeat(7, sig_892) and "0111010") or
		(repeat(7, sig_902) and "0100101") or
		(repeat(7, sig_899) and "0001101") or
		(repeat(7, sig_888) and "0110001") or
		(repeat(7, sig_886) and "0011011") or
		(repeat(7, sig_884) and "1001110") or
		(repeat(7, sig_878) and "0111101") or
		(repeat(7, sig_877) and "0101010") or
		(repeat(7, sig_876) and "0001001");

	-- Behaviour of component 'mux_377' model 'mux'
	mux_377 <=
		(repeat(32, sig_903) and decode_xa1_100(45 downto 14)) or
		(repeat(32, sig_1087) and decode_xa2_101(45 downto 14));

	-- Behaviour of component 'mux_372' model 'mux'
	mux_372 <=
		(repeat(32, sig_1081) and "00000000000000000000000001100100") or
		(repeat(32, sig_1087) and sig_1289(30 downto 0) & augh_main_i_132(0)) or
		(repeat(32, sig_950) and sig_1298(30 downto 0) & augh_main_i_132(0)) or
		(repeat(32, sig_1023) and sig_1288(30 downto 0) & augh_main_i_132(0));

	-- Behaviour of component 'mux_374' model 'mux'
	mux_374 <=
		(repeat(7, sig_903) and augh_main_i_132(6 downto 0)) or
		(repeat(7, sig_1087) and sig_1298(6 downto 0));

	-- Behaviour of component 'mux_364' model 'mux'
	mux_364 <=
		(repeat(32, sig_925) and "00000000000000000000000001111111") or
		(repeat(32, sig_914) and dec_del_dltx_reg1) or
		(repeat(32, sig_1253) and "00000000000000000000000000000000") or
		(repeat(32, sig_1016) and "00000000000000000000000000000000") or
		(repeat(32, sig_1241) and delay_dltx_reg1) or
		(repeat(32, sig_1195) and "00000000000000000000000000000000") or
		(repeat(32, sig_1129) and "00000000000000000000000011111111") or
		(repeat(32, sig_1133) and dec_del_dhx_reg1) or
		(repeat(32, sig_1153) and "00000000000000000000001000110100") or
		(repeat(32, sig_895) and dec_del_dhx_reg0) or
		(repeat(32, sig_868) and delay_dltx_reg0);

	-- Behaviour of component 'mux_365' model 'mux'
	mux_365 <=
		(repeat(33, sig_1112) and delay_bph_reg2(31) & delay_bph_reg2) or
		(repeat(33, sig_1125) and delay_bpl_reg2(31) & delay_bpl_reg2) or
		(repeat(33, sig_1153) and plt(31) & plt) or
		(repeat(33, sig_895) and dec_nbh(31) & dec_nbh) or
		(repeat(33, sig_932) and dec_del_bph_reg5(31) & dec_del_bph_reg5) or
		(repeat(33, sig_1053) and dec_del_bpl_reg5(31) & dec_del_bpl_reg5);

	-- Behaviour of component 'mux_366' model 'mux'
	mux_366 <=
		(repeat(32, sig_895) and "00000000000000000000000001111111") or
		(repeat(32, sig_1129) and "00000000000000000000000011111111") or
		(repeat(32, sig_1153) and plt2);

	-- Behaviour of component 'mux_363' model 'mux'
	mux_363 <=
		(repeat(33, sig_1016) and delay_bpl_reg4(31) & delay_bpl_reg4) or
		(repeat(33, sig_932) and dec_del_bph_reg3(31) & dec_del_bph_reg3) or
		(repeat(33, sig_1253) and delay_bpl_reg5(31) & delay_bpl_reg5) or
		(repeat(33, sig_1053) and dec_del_bpl_reg3(31) & dec_del_bpl_reg3) or
		(repeat(33, sig_1240) and delay_bpl_reg1(31) & delay_bpl_reg1) or
		(repeat(33, sig_1195) and delay_bpl_reg3(31) & delay_bpl_reg3) or
		(repeat(33, sig_1112) and delay_bph_reg1(31) & delay_bph_reg1) or
		(repeat(33, sig_1133) and dec_del_bph_reg1(31) & dec_del_bph_reg1) or
		(repeat(33, sig_1153) and deth(31) & deth) or
		(repeat(33, sig_927) and al2(31) & al2) or
		(repeat(33, sig_914) and dec_del_bpl_reg1(31) & dec_del_bpl_reg1) or
		(repeat(33, sig_911) and dec_nbl(31) & dec_nbl) or
		(repeat(33, sig_895) and dec_del_bph_reg0(31) & dec_del_bph_reg0) or
		(repeat(33, sig_868) and delay_bpl_reg0(31) & delay_bpl_reg0) or
		(repeat(33, sig_866) and delay_bpl_reg2(31) & delay_bpl_reg2);

	-- Behaviour of component 'mux_352' model 'mux'
	mux_352 <=
		(repeat(64, sig_1023) and "0000000000000000000000000000000000000000000000000000000000000001") or
		(repeat(64, sig_1133) and "0000000000000000000000000000000000000000000000000000000000000011") or
		(repeat(64, sig_1227) and sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31 downto 0)) or
		(repeat(64, sig_921) and filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45 downto 14)) or
		(repeat(64, sig_927) and sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38) & sig_1291(38 downto 7)) or
		(repeat(64, sig_954) and rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh(31) & rh);

	-- Behaviour of component 'mux_353' model 'mux'
	mux_353 <=
		(repeat(64, sig_926) and filtep_pl_14) or
		(repeat(64, sig_905) and dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt(31) & dec_dlt) or
		(repeat(64, sig_1145) and decode_xa2_101) or
		(repeat(64, sig_1022) and uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31 downto 6)) or
		(repeat(64, sig_1260) and encode_xb_68) or
		(repeat(64, sig_1198) and encode_xa_67) or
		(repeat(64, sig_1066) and decode_xa1_100) or
		(repeat(64, sig_1087) and augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31 downto 1)) or
		(repeat(64, sig_1133) and logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58(31) & logsch_wd_58) or
		(repeat(64, sig_893) and filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46 downto 15));

	-- Behaviour of component 'mux_354' model 'mux'
	mux_354 <=
		(repeat(64, sig_1087) and "0000000000000000000000000000000000000000000000000000000000000001") or
		(repeat(64, sig_1133) and sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308(31) & sig_1308) or
		(repeat(64, sig_1197) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31 downto 0)) or
		(repeat(64, sig_910) and filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45) & filtez_zl(45 downto 14)) or
		(repeat(64, sig_926) and sig_1303) or
		(repeat(64, sig_1022) and "0000000000000000000000000000000000000000000000000000000000000011");

	-- Behaviour of component 'mux_355' model 'mux'
	mux_355 <=
		(repeat(64, sig_927) and uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31 downto 6)) or
		(repeat(64, sig_1133) and filtez_zl) or
		(repeat(64, sig_1241) and filtep_pl_14);

	-- Behaviour of component 'mux_356' model 'mux'
	mux_356 <=
		(repeat(64, sig_927) and "0000000000000000000000000000000000000000000000000000000000000011") or
		(repeat(64, sig_1133) and sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31 downto 0)) or
		(repeat(64, sig_1241) and sig_1281);

	-- Behaviour of component 'mux_349' model 'mux'
	mux_349 <=
		(repeat(33, sig_1112) and delay_bph_reg3(31) & delay_bph_reg3) or
		(repeat(33, sig_1125) and delay_bpl_reg3(31) & delay_bpl_reg3) or
		(repeat(33, sig_1153) and nbh(31) & nbh) or
		(repeat(33, sig_895) and dec_rh1(30) & dec_rh1 & '0') or
		(repeat(33, sig_932) and dec_del_bph_reg2(31) & dec_del_bph_reg2) or
		(repeat(33, sig_1053) and dec_del_bpl_reg2(31) & dec_del_bpl_reg2);

	-- Behaviour of component 'mux_350' model 'mux'
	mux_350 <=
		(repeat(32, sig_895) and dec_ah1) or
		(repeat(32, sig_1129) and "00000000000000000000000011111111") or
		(repeat(32, sig_1153) and "00000000000000000000000001111111");

	-- Behaviour of component 'mux_351' model 'mux'
	mux_351 <=
		(repeat(64, sig_1023) and augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31) & augh_main_i_132(31 downto 1)) or
		(repeat(64, sig_1133) and uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31) & uppol1_wd2_51(31 downto 6)) or
		(repeat(64, sig_1227) and filtez_zl) or
		(repeat(64, sig_921) and filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46) & filtep_pl_14(46 downto 15)) or
		(repeat(64, sig_927) and uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42(31) & uppol2_wd4_42) or
		(repeat(64, sig_954) and rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl(31) & rl);

	-- Behaviour of component 'mux_341' model 'mux'
	mux_341 <=
		(repeat(64, sig_1045) and abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3) or
		(repeat(64, sig_1094) and uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53(31) & uppol1_apl1_53) or
		(repeat(64, sig_1142) and uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43) or
		(repeat(64, sig_1015) and "0000000000000000000000000000000000000000000000000000000000001010");

	-- Behaviour of component 'mux_342' model 'mux'
	mux_342 <=
		(repeat(64, sig_1045) and encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69(31) & encode_decis_69) or
		(repeat(64, sig_1094) and sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31) & sig_1307(31 downto 0)) or
		(repeat(64, sig_1142) and "1111111111111111111111111111111111111111111111111101000000000000") or
		(repeat(64, sig_1015) and sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5) & sig_1307(5 downto 0));

	-- Behaviour of component 'mux_338' model 'mux'
	mux_338 <=
		(repeat(32, sig_1257) and dec_dh);

	-- Behaviour of component 'mux_336' model 'mux'
	mux_336 <=
		(repeat(32, sig_1257) and dec_del_dhx_reg0);

	-- Behaviour of component 'mux_320' model 'mux'
	mux_320 <=
		(repeat(32, sig_932) and sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31 downto 8)) or
		(repeat(32, sig_1161) and sig_1298(31 downto 0));

	-- Behaviour of component 'mux_322' model 'mux'
	mux_322 <=
		(repeat(32, sig_932) and sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31 downto 8)) or
		(repeat(32, sig_974) and sig_1298(31 downto 0));

	-- Behaviour of component 'mux_324' model 'mux'
	mux_324 <=
		(repeat(32, sig_861) and sig_1298(31 downto 0)) or
		(repeat(32, sig_932) and sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31 downto 8));

	-- Behaviour of component 'mux_326' model 'mux'
	mux_326 <=
		(repeat(32, sig_862) and sig_1298(31 downto 0)) or
		(repeat(32, sig_932) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 8));

	-- Behaviour of component 'mux_310' model 'mux'
	mux_310 <=
		(repeat(32, sig_895) and dec_dlt);

	-- Behaviour of component 'mux_314' model 'mux'
	mux_314 <=
		(repeat(33, sig_927) and plt(31) & plt) or
		(repeat(33, sig_911) and dec_detl(31) & dec_detl) or
		(repeat(33, sig_1133) and dec_al2(31) & dec_al2) or
		(repeat(33, sig_932) and dec_del_bph_reg1(31) & dec_del_bph_reg1) or
		(repeat(33, sig_1153) and al1(31) & al1) or
		(repeat(33, sig_1241) and rlt2(30) & rlt2 & '0') or
		(repeat(33, sig_1053) and dec_del_bpl_reg1(31) & dec_del_bpl_reg1) or
		(repeat(33, sig_1112) and delay_bph_reg4(31) & delay_bph_reg4) or
		(repeat(33, sig_1125) and delay_bpl_reg4(31) & delay_bpl_reg4) or
		(repeat(33, sig_895) and dec_al1(31) & dec_al1) or
		(repeat(33, sig_868) and rlt1(30) & rlt1 & '0');

	-- Behaviour of component 'mux_315' model 'mux'
	mux_315 <=
		(repeat(32, sig_1133) and "00000000000000000000000001111111") or
		(repeat(32, sig_1150) and "00000000000000000000000011111111") or
		(repeat(32, sig_1241) and al2) or
		(repeat(32, sig_868) and al1) or
		(repeat(32, sig_911) and sig_1315) or
		(repeat(32, sig_927) and plt1);

	-- Behaviour of component 'mux_316' model 'mux'
	mux_316 <=
		(repeat(32, sig_932) and sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31 downto 8)) or
		(repeat(32, sig_1171) and sig_1298(31 downto 0));

	-- Behaviour of component 'mux_318' model 'mux'
	mux_318 <=
		(repeat(32, sig_890) and sig_1298(31 downto 0)) or
		(repeat(32, sig_932) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31 downto 8));

	-- Behaviour of component 'mux_308' model 'mux'
	mux_308 <=
		(repeat(32, sig_895) and dec_del_dltx_reg0);

	-- Behaviour of component 'mux_292' model 'mux'
	mux_292 <=
		(repeat(32, sig_1017) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1053) and sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31 downto 8));

	-- Behaviour of component 'mux_294' model 'mux'
	mux_294 <=
		(repeat(32, sig_1053) and sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31 downto 8)) or
		(repeat(32, sig_1268) and sig_1298(31 downto 0));

	-- Behaviour of component 'mux_296' model 'mux'
	mux_296 <=
		(repeat(32, sig_871) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1053) and sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31 downto 8));

	-- Behaviour of component 'mux_298' model 'mux'
	mux_298 <=
		(repeat(32, sig_1053) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 8)) or
		(repeat(32, sig_1262) and sig_1298(31 downto 0));

	-- Behaviour of component 'mux_290' model 'mux'
	mux_290 <=
		(repeat(32, sig_1053) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31 downto 8)) or
		(repeat(32, sig_1174) and sig_1298(31 downto 0));

	-- Behaviour of component 'mux_286' model 'mux'
	mux_286 <=
		(repeat(32, sig_864) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1112) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 8));

	-- Behaviour of component 'mux_288' model 'mux'
	mux_288 <=
		(repeat(32, sig_936) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1053) and sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31 downto 8));

	-- Behaviour of component 'mux_284' model 'mux'
	mux_284 <=
		(repeat(32, sig_1112) and sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31 downto 8)) or
		(repeat(32, sig_1280) and sig_1298(31 downto 0));

	-- Behaviour of component 'mux_278' model 'mux'
	mux_278 <=
		(repeat(32, sig_875) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1112) and sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31 downto 8));

	-- Behaviour of component 'mux_280' model 'mux'
	mux_280 <=
		(repeat(32, sig_1000) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1112) and sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31 downto 8));

	-- Behaviour of component 'mux_282' model 'mux'
	mux_282 <=
		(repeat(32, sig_863) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1112) and sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31 downto 8));

	-- Behaviour of component 'mux_272' model 'mux'
	mux_272 <=
		(repeat(32, sig_997) and delay_dhx_reg0);

	-- Behaviour of component 'mux_274' model 'mux'
	mux_274 <=
		(repeat(32, sig_997) and dh);

	-- Behaviour of component 'mux_276' model 'mux'
	mux_276 <=
		(repeat(32, sig_1092) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1112) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31 downto 8));

	-- Behaviour of component 'mux_262' model 'mux'
	mux_262 <=
		(repeat(32, sig_1153) and dlt);

	-- Behaviour of component 'mux_260' model 'mux'
	mux_260 <=
		(repeat(32, sig_1153) and delay_dltx_reg0);

	-- Behaviour of component 'mux_250' model 'mux'
	mux_250 <=
		(repeat(32, sig_923) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1125) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 8));

	-- Behaviour of component 'mux_248' model 'mux'
	mux_248 <=
		(repeat(32, sig_1042) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1125) and sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31 downto 8));

	-- Behaviour of component 'mux_244' model 'mux'
	mux_244 <=
		(repeat(32, sig_1036) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1125) and sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31) & sig_1287(31 downto 8));

	-- Behaviour of component 'mux_246' model 'mux'
	mux_246 <=
		(repeat(32, sig_1040) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1125) and sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31) & sig_1292(31 downto 8));

	-- Behaviour of component 'mux_242' model 'mux'
	mux_242 <=
		(repeat(32, sig_1086) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1125) and sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31 downto 8));

	-- Behaviour of component 'mux_238' model 'mux'
	mux_238 <=
		(repeat(32, sig_1008) and xd);

	-- Behaviour of component 'mux_240' model 'mux'
	mux_240 <=
		(repeat(32, sig_1199) and sig_1298(31 downto 0)) or
		(repeat(32, sig_1125) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31 downto 8));

	-- Behaviour of component 'mux_236' model 'mux'
	mux_236 <=
		(repeat(32, sig_1008) and accumc_reg0);

	-- Behaviour of component 'mux_232' model 'mux'
	mux_232 <=
		(repeat(32, sig_1008) and accumc_reg2);

	-- Behaviour of component 'mux_234' model 'mux'
	mux_234 <=
		(repeat(32, sig_1008) and accumc_reg1);

	-- Behaviour of component 'mux_230' model 'mux'
	mux_230 <=
		(repeat(32, sig_1008) and accumc_reg3);

	-- Behaviour of component 'mux_226' model 'mux'
	mux_226 <=
		(repeat(32, sig_1008) and accumc_reg5);

	-- Behaviour of component 'mux_228' model 'mux'
	mux_228 <=
		(repeat(32, sig_1008) and accumc_reg4);

	-- Behaviour of component 'mux_224' model 'mux'
	mux_224 <=
		(repeat(32, sig_1008) and accumc_reg6);

	-- Behaviour of component 'mux_220' model 'mux'
	mux_220 <=
		(repeat(32, sig_1008) and accumc_reg8);

	-- Behaviour of component 'mux_222' model 'mux'
	mux_222 <=
		(repeat(32, sig_1008) and accumc_reg7);

	-- Behaviour of component 'mux_218' model 'mux'
	mux_218 <=
		(repeat(32, sig_1008) and accumc_reg9);

	-- Behaviour of component 'mux_214' model 'mux'
	mux_214 <=
		(repeat(32, sig_1008) and accumd_reg0);

	-- Behaviour of component 'mux_216' model 'mux'
	mux_216 <=
		(repeat(32, sig_1008) and xs);

	-- Behaviour of component 'mux_212' model 'mux'
	mux_212 <=
		(repeat(32, sig_1008) and accumd_reg1);

	-- Behaviour of component 'mux_208' model 'mux'
	mux_208 <=
		(repeat(32, sig_1008) and accumd_reg3);

	-- Behaviour of component 'mux_210' model 'mux'
	mux_210 <=
		(repeat(32, sig_1008) and accumd_reg2);

	-- Behaviour of component 'mux_206' model 'mux'
	mux_206 <=
		(repeat(32, sig_1008) and accumd_reg4);

	-- Behaviour of component 'mux_202' model 'mux'
	mux_202 <=
		(repeat(32, sig_1008) and accumd_reg6);

	-- Behaviour of component 'mux_204' model 'mux'
	mux_204 <=
		(repeat(32, sig_1008) and accumd_reg5);

	-- Behaviour of component 'mux_200' model 'mux'
	mux_200 <=
		(repeat(32, sig_1008) and accumd_reg7);

	-- Behaviour of component 'mux_196' model 'mux'
	mux_196 <=
		(repeat(32, sig_1008) and accumd_reg9);

	-- Behaviour of component 'mux_198' model 'mux'
	mux_198 <=
		(repeat(32, sig_1008) and accumd_reg8);

	-- Behaviour of component 'mux_194' model 'mux'
	mux_194 <=
		(repeat(32, sig_1175) and tqmf_reg6);

	-- Behaviour of component 'mux_190' model 'mux'
	mux_190 <=
		(repeat(32, sig_1175) and tqmf_reg8);

	-- Behaviour of component 'mux_192' model 'mux'
	mux_192 <=
		(repeat(32, sig_1175) and tqmf_reg7);

	-- Behaviour of component 'mux_188' model 'mux'
	mux_188 <=
		(repeat(32, sig_1175) and tqmf_reg9);

	-- Behaviour of component 'mux_184' model 'mux'
	mux_184 <=
		(repeat(32, sig_1175) and tqmf_reg11);

	-- Behaviour of component 'mux_186' model 'mux'
	mux_186 <=
		(repeat(32, sig_1175) and tqmf_reg10);

	-- Behaviour of component 'mux_182' model 'mux'
	mux_182 <=
		(repeat(32, sig_1175) and tqmf_reg12);

	-- Behaviour of component 'mux_178' model 'mux'
	mux_178 <=
		(repeat(32, sig_1175) and tqmf_reg14);

	-- Behaviour of component 'mux_180' model 'mux'
	mux_180 <=
		(repeat(32, sig_1175) and tqmf_reg13);

	-- Behaviour of component 'mux_176' model 'mux'
	mux_176 <=
		(repeat(32, sig_1175) and tqmf_reg15);

	-- Behaviour of component 'mux_172' model 'mux'
	mux_172 <=
		(repeat(32, sig_1175) and tqmf_reg17);

	-- Behaviour of component 'mux_174' model 'mux'
	mux_174 <=
		(repeat(32, sig_1175) and tqmf_reg16);

	-- Behaviour of component 'mux_170' model 'mux'
	mux_170 <=
		(repeat(32, sig_1175) and tqmf_reg18);

	-- Behaviour of component 'mux_166' model 'mux'
	mux_166 <=
		(repeat(32, sig_1175) and tqmf_reg20);

	-- Behaviour of component 'mux_168' model 'mux'
	mux_168 <=
		(repeat(32, sig_1175) and tqmf_reg19);

	-- Behaviour of component 'mux_164' model 'mux'
	mux_164 <=
		(repeat(32, sig_1175) and tqmf_reg21);

	-- Behaviour of component 'not_709' model 'not'
	not_709 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'or_710' model 'or'
	or_710 <=
		and_713 or
		and_711;

	-- Behaviour of component 'or_692' model 'or'
	or_692 <=
		sig_1303(31) & "0000000" or
		not_693 & "0000000";

	-- Behaviour of component 'not_693' model 'not'
	not_693 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'not_768' model 'not'
	not_768 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'or_769' model 'or'
	or_769 <=
		and_771 or
		and_770;

	-- Behaviour of component 'and_770' model 'and'
	and_770 <=
		uppol1_wd3_52 and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'and_771' model 'and'
	and_771 <=
		uppol1_apl1_53 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'or_619' model 'or'
	or_619 <=
		sig_1303(31) & "0000000" or
		not_620 & "0000000";

	-- Behaviour of component 'not_620' model 'not'
	not_620 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'or_621' model 'or'
	or_621 <=
		sig_1304(31) & "0000000" or
		not_622 & "0000000";

	-- Behaviour of component 'not_622' model 'not'
	not_622 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'or_623' model 'or'
	or_623 <=
		sig_1303(31) & "0000000" or
		not_624 & "0000000";

	-- Behaviour of component 'not_624' model 'not'
	not_624 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'or_625' model 'or'
	or_625 <=
		sig_1304(31) & "0000000" or
		not_626 & "0000000";

	-- Behaviour of component 'not_626' model 'not'
	not_626 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'or_627' model 'or'
	or_627 <=
		sig_1304(31) & "0000000" or
		not_628 & "0000000";

	-- Behaviour of component 'and_633' model 'and'
	and_633 <=
		uppol2_apl2_43 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'not_628' model 'not'
	not_628 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'or_629' model 'or'
	or_629 <=
		sig_1304(31) & "0000000" or
		not_630 & "0000000";

	-- Behaviour of component 'not_630' model 'not'
	not_630 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'or_631' model 'or'
	or_631 <=
		and_633 or
		and_632;

	-- Behaviour of component 'or_634' model 'or'
	or_634 <=
		sig_1304(31) & "0000000" or
		not_635 & "0000000";

	-- Behaviour of component 'not_635' model 'not'
	not_635 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'or_636' model 'or'
	or_636 <=
		sig_1292(31) & "0000000" or
		not_637 & "0000000";

	-- Behaviour of component 'not_637' model 'not'
	not_637 <= not (
		sig_1292(31)
	);

	-- Behaviour of component 'and_632' model 'and'
	and_632 <=
		"00000000000000000011000000000000" and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'or_641' model 'or'
	or_641 <=
		and_643 or
		and_642;

	-- Behaviour of component 'and_640' model 'and'
	and_640 <=
		logsch_nbh_57 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'and_645' model 'and'
	and_645 <=
		sig_1288(25 downto 0) & uppol1_wd2_51(5 downto 0) and
		not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646 & not_646;

	-- Behaviour of component 'and_639' model 'and'
	and_639 <=
		"00000000000000000101100000000000" and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'and_643' model 'and'
	and_643 <=
		uppol2_apl2_43 and
		sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317 & sig_1317;

	-- Behaviour of component 'and_650' model 'and'
	and_650 <=
		logscl_nbl_27 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'or_651' model 'or'
	or_651 <=
		and_653 or
		and_652;

	-- Behaviour of component 'or_644' model 'or'
	or_644 <=
		and_647 or
		and_645;

	-- Behaviour of component 'and_649' model 'and'
	and_649 <=
		"00000000000000000100100000000000" and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'mux_498' model 'mux'
	mux_498 <=
		(repeat(32, sig_1133) and dec_plt);

	-- Behaviour of component 'mux_500' model 'mux'
	mux_500 <=
		(repeat(32, sig_895) and dec_plt1);

	-- Behaviour of component 'mux_502' model 'mux'
	mux_502 <=
		(repeat(32, sig_990) and "00000000000000000000000000001000") or
		(repeat(32, sig_1101) and scalel_wd3_35 & "000");

	-- Behaviour of component 'mux_504' model 'mux'
	mux_504 <=
		(repeat(32, sig_990) and "00000000000000000000000000100000") or
		(repeat(32, sig_1122) and scalel_wd3_35 & "000");

	-- Behaviour of component 'and_652' model 'and'
	and_652 <=
		uppol1_wd3_52 and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'and_653' model 'and'
	and_653 <=
		uppol1_apl1_53 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'or_654' model 'or'
	or_654 <=
		and_656 or
		and_655;

	-- Behaviour of component 'and_655' model 'and'
	and_655 <=
		sig_1307(31 downto 0) and
		sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301;

	-- Behaviour of component 'and_656' model 'and'
	and_656 <=
		uppol1_apl1_53 and
		sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282;

	-- Behaviour of component 'or_657' model 'or'
	or_657 <=
		and_659 or
		and_658;

	-- Behaviour of component 'and_658' model 'and'
	and_658 <=
		"00000000000000000011000000000000" and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'and_659' model 'and'
	and_659 <=
		uppol2_apl2_43 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'mux_510' model 'mux'
	mux_510 <=
		(repeat(31, sig_1023) and yh);

	-- Behaviour of component 'mux_512' model 'mux'
	mux_512 <=
		(repeat(31, sig_997) and rh1);

	-- Behaviour of component 'not_661' model 'not'
	not_661 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'and_665' model 'and'
	and_665 <=
		uppol1_apl1_53 and
		sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282;

	-- Behaviour of component 'or_666' model 'or'
	or_666 <=
		and_668 or
		and_667;

	-- Behaviour of component 'mux_514' model 'mux'
	mux_514 <=
		(repeat(32, sig_1023) and ph);

	-- Behaviour of component 'mux_516' model 'mux'
	mux_516 <=
		(repeat(32, sig_997) and ph1);

	-- Behaviour of component 'mux_518' model 'mux'
	mux_518 <=
		(repeat(32, sig_995) and uppol1_apl1_53);

	-- Behaviour of component 'mux_520' model 'mux'
	mux_520 <=
		(repeat(32, sig_1005) and uppol2_apl2_43);

	-- Behaviour of component 'and_647' model 'and'
	and_647 <=
		sig_1302(31 downto 0) and
		sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31);

	-- Behaviour of component 'and_664' model 'and'
	and_664 <=
		sig_1307(31 downto 0) and
		sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301;

	-- Behaviour of component 'and_667' model 'and'
	and_667 <=
		"00000000000000000101100000000000" and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'and_670' model 'and'
	and_670 <=
		sig_1311 and
		not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671 & not_671;

	-- Behaviour of component 'and_672' model 'and'
	and_672 <=
		sig_1310 and
		quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16 & quantl_el_16;

	-- Behaviour of component 'or_674' model 'or'
	or_674 <=
		and_676 or
		and_675;

	-- Behaviour of component 'mux_528' model 'mux'
	mux_528 <=
		(repeat(32, sig_1069) and logsch_nbh_57);

	-- Behaviour of component 'or_638' model 'or'
	or_638 <=
		and_640 or
		and_639;

	-- Behaviour of component 'and_642' model 'and'
	and_642 <=
		"11111111111111111101000000000000" and
		sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284 & sig_1284;

	-- Behaviour of component 'or_648' model 'or'
	or_648 <=
		and_650 or
		and_649;

	-- Behaviour of component 'or_669' model 'or'
	or_669 <=
		and_672 or
		and_670;

	-- Behaviour of component 'and_676' model 'and'
	and_676 <=
		ih and
		sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283 & sig_1283;

	-- Behaviour of component 'mux_532' model 'mux'
	mux_532 <=
		(repeat(32, sig_914) and decode_input_98(29) & decode_input_98(29) & decode_input_98(29) & decode_input_98(29) & decode_input_98(29) & decode_input_98(29) & decode_input_98(29 downto 4)) or
		(repeat(32, sig_976) and or_701) or
		(repeat(32, sig_1045) and or_674);

	-- Behaviour of component 'mux_534' model 'mux'
	mux_534 <=
		(repeat(2, sig_869) and ih(1 downto 0)) or
		(repeat(2, sig_1133) and decode_input_98(5 downto 4));

	-- Behaviour of component 'mux_535' model 'mux'
	mux_535 <=
		(repeat(2, sig_869) and ih(1 downto 0)) or
		(repeat(2, sig_895) and decode_input_98(5 downto 4));

	-- Behaviour of component 'or_663' model 'or'
	or_663 <=
		and_665 or
		and_664;

	-- Behaviour of component 'and_668' model 'and'
	and_668 <=
		logsch_nbh_57 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'or_679' model 'or'
	or_679 <=
		sig_1304(31) & "0000000" or
		not_680 & "0000000";

	-- Behaviour of component 'not_680' model 'not'
	not_680 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'not_682' model 'not'
	not_682 <= not (
		logscl_nbl_27(31)
	);

	-- Behaviour of component 'or_683' model 'or'
	or_683 <=
		sig_1303(31) & "0000000" or
		not_684 & "0000000";

	-- Behaviour of component 'and_686' model 'and'
	and_686 <=
		"00000000000000000100100000000000" and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'and_689' model 'and'
	and_689 <=
		sig_1289(25 downto 0) & uppol1_wd2_51(5 downto 0) and
		not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690 & not_690;

	-- Behaviour of component 'mux_540' model 'mux'
	mux_540 <=
		(repeat(32, sig_990) and "00000000000000000000000000001000") or
		(repeat(32, sig_1057) and scalel_wd3_35 & "000");

	-- Behaviour of component 'mux_544' model 'mux'
	mux_544 <=
		(repeat(32, sig_990) and "00000000000000000000000000100000") or
		(repeat(32, sig_1011) and scalel_wd3_35 & "000");

	-- Behaviour of component 'or_660' model 'or'
	or_660 <=
		sig_1303(31) & "0000000" or
		not_661 & "0000000";

	-- Behaviour of component 'or_677' model 'or'
	or_677 <=
		sig_1304(31) & "0000000" or
		not_678 & "0000000";

	-- Behaviour of component 'not_678' model 'not'
	not_678 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'not_684' model 'not'
	not_684 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'or_685' model 'or'
	or_685 <=
		and_687 or
		and_686;

	-- Behaviour of component 'or_688' model 'or'
	or_688 <=
		and_691 or
		and_689;

	-- Behaviour of component 'or_695' model 'or'
	or_695 <=
		sig_1303(31) & "0000000" or
		not_696 & "0000000";

	-- Behaviour of component 'not_671' model 'not'
	not_671 <= not (
		quantl_el_16
	);

	-- Behaviour of component 'not_696' model 'not'
	not_696 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'or_697' model 'or'
	or_697 <=
		sig_1304(31) & "0000000" or
		not_698 & "0000000";

	-- Behaviour of component 'not_698' model 'not'
	not_698 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'or_699' model 'or'
	or_699 <=
		ih(25 downto 0) or
		quantl_ril_18(31 downto 6);

	-- Behaviour of component 'not_703' model 'not'
	not_703 <= not (
		eh(31)
	);

	-- Behaviour of component 'mux_563' model 'mux'
	mux_563 <=
		(repeat(32, sig_1003) and uppol2_apl2_43);

	-- Behaviour of component 'mux_549' model 'mux'
	mux_549 <=
		(repeat(31, sig_927) and rlt);

	-- Behaviour of component 'mux_551' model 'mux'
	mux_551 <=
		(repeat(31, sig_1153) and rlt1);

	-- Behaviour of component 'mux_557' model 'mux'
	mux_557 <=
		(repeat(32, sig_927) and plt);

	-- Behaviour of component 'mux_559' model 'mux'
	mux_559 <=
		(repeat(32, sig_1153) and plt1);

	-- Behaviour of component 'mux_561' model 'mux'
	mux_561 <=
		(repeat(32, sig_964) and uppol1_apl1_53);

	-- Behaviour of component 'not_646' model 'not'
	not_646 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'and_675' model 'and'
	and_675 <=
		sig_1307(31 downto 0) and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'and_681' model 'and'
	and_681 <=
		logscl_nbl_27 and
		not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682 & not_682;

	-- Behaviour of component 'not_690' model 'not'
	not_690 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'and_691' model 'and'
	and_691 <=
		sig_1302(31 downto 0) and
		sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31);

	-- Behaviour of component 'and_702' model 'and'
	and_702 <=
		"00000000000000000000000000000011" and
		not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703;

	-- Behaviour of component 'or_705' model 'or'
	or_705 <=
		and_707 or
		and_706;

	-- Behaviour of component 'not_712' model 'not'
	not_712 <= not (
		el(31)
	);

	-- Behaviour of component 'or_717' model 'or'
	or_717 <=
		and_719 or
		and_718;

	-- Behaviour of component 'not_722' model 'not'
	not_722 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'mux_565' model 'mux'
	mux_565 <=
		(repeat(32, sig_891) and logscl_nbl_27);

	-- Behaviour of component 'mux_567' model 'mux'
	mux_567 <=
		(repeat(5, sig_1031) and logscl_nbl_27(10 downto 6)) or
		(repeat(5, sig_1070) and logsch_nbh_57(10 downto 6));

	-- Behaviour of component 'mux_568' model 'mux'
	mux_568 <=
		(repeat(4, sig_914) and decode_input_98(3 downto 0)) or
		(repeat(4, sig_1100) and quantl_ril_18(5 downto 2));

	-- Behaviour of component 'mux_570' model 'mux'
	mux_570 <=
		(repeat(4, sig_914) and decode_input_98(3 downto 0)) or
		(repeat(4, sig_1100) and quantl_ril_18(5 downto 2));

	-- Behaviour of component 'and_687' model 'and'
	and_687 <=
		logscl_nbl_27 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'and_704' model 'and'
	and_704 <=
		"00000000000000000000000000000001" and
		eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31);

	-- Behaviour of component 'and_707' model 'and'
	and_707 <=
		sig_1302(31 downto 0) and
		eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31) & eh(31);

	-- Behaviour of component 'and_716' model 'and'
	and_716 <=
		uppol2_apl2_43 and
		sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305;

	-- Behaviour of component 'or_720' model 'or'
	or_720 <=
		and_723 or
		and_721;

	-- Behaviour of component 'and_721' model 'and'
	and_721 <=
		sig_1289(25 downto 0) & uppol1_wd2_51(5 downto 0) and
		not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722 & not_722;

	-- Behaviour of component 'and_724' model 'and'
	and_724 <=
		logscl_nbl_27 and
		not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725 & not_725;

	-- Behaviour of component 'or_730' model 'or'
	or_730 <=
		sig_1304(31) & "0000000" or
		not_731 & "0000000";

	-- Behaviour of component 'not_731' model 'not'
	not_731 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'or_732' model 'or'
	or_732 <=
		sig_1304(31) & "0000000" or
		not_733 & "0000000";

	-- Behaviour of component 'not_733' model 'not'
	not_733 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'or_734' model 'or'
	or_734 <=
		and_736 or
		and_735;

	-- Behaviour of component 'or_740' model 'or'
	or_740 <=
		sig_1303(31) & "0000000" or
		not_741 & "0000000";

	-- Behaviour of component 'not_741' model 'not'
	not_741 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'and_706' model 'and'
	and_706 <=
		eh and
		not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703 & not_703;

	-- Behaviour of component 'and_713' model 'and'
	and_713 <=
		sig_1302(31 downto 0) and
		el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31) & el(31);

	-- Behaviour of component 'and_718' model 'and'
	and_718 <=
		"00000000000000000011000000000000" and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'and_719' model 'and'
	and_719 <=
		uppol2_apl2_43 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'not_725' model 'not'
	not_725 <= not (
		logscl_nbl_27(31)
	);

	-- Behaviour of component 'or_726' model 'or'
	or_726 <=
		and_729 or
		and_727;

	-- Behaviour of component 'mux_587' model 'mux'
	mux_587 <=
		(repeat(32, sig_1042) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_677) or
		(repeat(32, sig_1040) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_679) or
		(repeat(32, sig_1268) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_623) or
		(repeat(32, sig_1086) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_660) or
		(repeat(32, sig_1270) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_621) or
		(repeat(32, sig_1280) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_619) or
		(repeat(32, sig_1161) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_634) or
		(repeat(32, sig_1174) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_629) or
		(repeat(32, sig_1262) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_625) or
		(repeat(32, sig_1036) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_683) or
		(repeat(32, sig_1017) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_692) or
		(repeat(32, sig_1000) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_695) or
		(repeat(32, sig_974) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_708) or
		(repeat(32, sig_923) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_730) or
		(repeat(32, sig_922) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_732) or
		(repeat(32, sig_890) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_745) or
		(repeat(32, sig_875) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_761) or
		(repeat(32, sig_872) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_765) or
		(repeat(32, sig_871) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_767) or
		(repeat(32, sig_864) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_772) or
		(repeat(32, sig_863) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_774) or
		(repeat(32, sig_862) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & or_776) or
		(repeat(32, sig_861) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_778) or
		(repeat(32, sig_1200) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & or_780);

	-- Behaviour of component 'mux_589' model 'mux'
	mux_589 <=
		(repeat(32, sig_1269) and sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31) & sig_1303(31 downto 8)) or
		(repeat(32, sig_1276) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 8));

	-- Behaviour of component 'mux_591' model 'mux'
	mux_591 <=
		(repeat(64, sig_1154) and sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 0)) or
		(repeat(64, sig_1169) and sig_1298) or
		(repeat(64, sig_1227) and sig_1288) or
		(repeat(64, sig_896) and sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31 downto 0)) or
		(repeat(64, sig_1133) and sig_1290);

	-- Behaviour of component 'mux_593' model 'mux'
	mux_593 <=
		(repeat(32, sig_949) and sig_1294) or
		(repeat(32, sig_1209) and sig_1293);

	-- Behaviour of component 'mux_597' model 'mux'
	mux_597 <=
		(repeat(32, sig_1175) and tqmf_reg5);

	-- Behaviour of component 'mux_599' model 'mux'
	mux_599 <=
		(repeat(32, sig_1175) and tqmf_reg4);

	-- Behaviour of component 'mux_601' model 'mux'
	mux_601 <=
		(repeat(32, sig_1175) and tqmf_reg3);

	-- Behaviour of component 'mux_603' model 'mux'
	mux_603 <=
		(repeat(32, sig_1175) and tqmf_reg2);

	-- Behaviour of component 'mux_605' model 'mux'
	mux_605 <=
		(repeat(32, sig_1175) and tqmf_reg1);

	-- Behaviour of component 'mux_607' model 'mux'
	mux_607 <=
		(repeat(32, sig_1175) and tqmf_reg0);

	-- Behaviour of component 'mux_609' model 'mux'
	mux_609 <=
		(repeat(32, sig_1175) and encode_xin1_61);

	-- Behaviour of component 'mux_611' model 'mux'
	mux_611 <=
		(repeat(32, sig_1175) and encode_xin2_62);

	-- Behaviour of component 'or_701' model 'or'
	or_701 <=
		and_704 or
		and_702;

	-- Behaviour of component 'or_708' model 'or'
	or_708 <=
		sig_1303(31) & "0000000" or
		not_709 & "0000000";

	-- Behaviour of component 'and_711' model 'and'
	and_711 <=
		el and
		not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712 & not_712;

	-- Behaviour of component 'and_729' model 'and'
	and_729 <=
		sig_1302(31 downto 0) and
		sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31);

	-- Behaviour of component 'and_736' model 'and'
	and_736 <=
		uppol1_apl1_53 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'or_737' model 'or'
	or_737 <=
		and_739 or
		and_738;

	-- Behaviour of component 'and_738' model 'and'
	and_738 <=
		"11111111111111111101000000000000" and
		sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301;

	-- Behaviour of component 'and_739' model 'and'
	and_739 <=
		uppol2_apl2_43 and
		sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305 & sig_1305;

	-- Behaviour of component 'or_745' model 'or'
	or_745 <=
		sig_1303(31) & "0000000" or
		not_746 & "0000000";

	-- Behaviour of component 'and_749' model 'and'
	and_749 <=
		uppol2_apl2_43 and
		sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306 & sig_1306;

	-- Behaviour of component 'and_750' model 'and'
	and_750 <=
		logsch_nbh_57 and
		not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751 & not_751;

	-- Behaviour of component 'and_754' model 'and'
	and_754 <=
		uppol1_apl1_53 and
		sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282 & sig_1282;

	-- Behaviour of component 'and_756' model 'and'
	and_756 <=
		uppol1_wd3_52 and
		sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299 & sig_1299;

	-- Behaviour of component 'and_759' model 'and'
	and_759 <=
		"11111111111111111101000000000000" and
		sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301 & sig_1301;

	-- Behaviour of component 'and_763' model 'and'
	and_763 <=
		logsch_nbh_57 and
		not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764 & not_764;

	-- Behaviour of component 'or_765' model 'or'
	or_765 <=
		sig_1304(31) & "0000000" or
		not_766 & "0000000";

	-- Behaviour of component 'or_772' model 'or'
	or_772 <=
		sig_1304(31) & "0000000" or
		not_773 & "0000000";

	-- Behaviour of component 'not_773' model 'not'
	not_773 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'or_774' model 'or'
	or_774 <=
		sig_1303(31) & "0000000" or
		not_775 & "0000000";

	-- Behaviour of component 'not_775' model 'not'
	not_775 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'or_776' model 'or'
	or_776 <=
		sig_1303(31) & "0000000" or
		not_777 & "0000000";

	-- Behaviour of component 'not_777' model 'not'
	not_777 <= not (
		sig_1303(31)
	);

	-- Behaviour of component 'or_778' model 'or'
	or_778 <=
		sig_1304(31) & "0000000" or
		not_779 & "0000000";

	-- Behaviour of component 'not_779' model 'not'
	not_779 <= not (
		sig_1304(31)
	);

	-- Behaviour of component 'or_780' model 'or'
	or_780 <=
		sig_1304(31) & "0000000" or
		not_781 & "0000000";

	-- Behaviour of component 'not_781' model 'not'
	not_781 <= not (
		sig_1304(31)
	);

	-- Behaviour of all components of model 'reg'
	-- Registers with clock = sig_clock and no reset
	process(sig_clock)
	begin
		if rising_edge(sig_clock) then
			if sig_1176 = '1' then
				tqmf_reg0 <= mux_611;
			end if;
			if sig_1176 = '1' then
				tqmf_reg1 <= mux_609;
			end if;
			if sig_1176 = '1' then
				tqmf_reg2 <= mux_607;
			end if;
			if sig_1176 = '1' then
				tqmf_reg3 <= mux_605;
			end if;
			if sig_1176 = '1' then
				tqmf_reg4 <= mux_603;
			end if;
			if sig_1176 = '1' then
				tqmf_reg5 <= mux_601;
			end if;
			if sig_1176 = '1' then
				tqmf_reg6 <= mux_599;
			end if;
			if sig_1176 = '1' then
				tqmf_reg7 <= mux_597;
			end if;
			if sig_1221 = '1' then
				read32_buf_0 <= stdin_data;
			end if;
			if sig_1215 = '1' then
				write32_val_1 <= mux_593;
			end if;
			if sig_1226 = '1' then
				filtez_zl <= mux_591;
			end if;
			if sig_1274 = '1' then
				upzero_wd3 <= mux_589;
			end if;
			if sig_1274 = '1' then
				upzero_wd2 <= mux_587;
			end if;
			if sig_956 = '1' then
				xh <= sig_1302(46 downto 15);
			end if;
			if sig_956 = '1' then
				xl <= sig_1298(46 downto 15);
			end if;
			if sig_953 = '1' then
				xd <= sig_1307(31 downto 0);
			end if;
			if sig_953 = '1' then
				xs <= sig_1288(31 downto 0);
			end if;
			if sig_958 = '1' then
				el <= sig_1302(31 downto 0);
			end if;
			if sig_920 = '1' then
				sl <= sig_1288(31 downto 0);
			end if;
			if sig_920 = '1' then
				szl <= filtez_zl(45 downto 14);
			end if;
			if sig_1098 = '1' then
				il <= quantl_ril_18(5 downto 0);
			end if;
			if sig_983 = '1' then
				nbl <= mux_565;
			end if;
			if sig_1001 = '1' then
				al2 <= mux_563;
			end if;
			if sig_984 = '1' then
				al1 <= mux_561;
			end if;
			if sig_1151 = '1' then
				plt2 <= mux_559;
			end if;
			if sig_989 = '1' then
				plt1 <= mux_557;
			end if;
			if sig_934 = '1' then
				plt <= sig_1298(31 downto 0);
			end if;
			if sig_1098 = '1' then
				dlt <= sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 15);
			end if;
			if sig_1151 = '1' then
				rlt2 <= mux_551;
			end if;
			if sig_989 = '1' then
				rlt1 <= mux_549;
			end if;
			if sig_1152 = '1' then
				rlt <= sig_1298(30 downto 0);
			end if;
			if sig_1010 = '1' then
				detl <= mux_544;
			end if;
			if sig_1056 = '1' then
				deth <= mux_540;
			end if;
			if sig_1095 = '1' then
				sh <= sig_1298(31 downto 0);
			end if;
			if sig_963 = '1' then
				eh <= sig_1302(31 downto 0);
			end if;
			if sig_1043 = '1' then
				ih <= mux_532;
			end if;
			if sig_870 = '1' then
				dh <= sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 15);
			end if;
			if sig_1071 = '1' then
				nbh <= mux_528;
			end if;
			if sig_1255 = '1' then
				rh <= sig_1298(31 downto 0);
			end if;
			if sig_996 = '1' then
				yh <= sig_1298(30 downto 0);
			end if;
			if sig_873 = '1' then
				ph <= sig_1298(31 downto 0);
			end if;
			if sig_1004 = '1' then
				ah2 <= mux_520;
			end if;
			if sig_994 = '1' then
				ah1 <= mux_518;
			end if;
			if sig_998 = '1' then
				ph2 <= mux_516;
			end if;
			if sig_1021 = '1' then
				ph1 <= mux_514;
			end if;
			if sig_998 = '1' then
				rh2 <= mux_512;
			end if;
			if sig_1021 = '1' then
				rh1 <= mux_510;
			end if;
			if sig_1083 = '1' then
				rl <= sig_1298(31 downto 0);
			end if;
			if sig_915 = '1' then
				dec_dlt <= sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 15);
			end if;
			if sig_1121 = '1' then
				dec_detl <= mux_504;
			end if;
			if sig_1105 = '1' then
				dec_deth <= mux_502;
			end if;
			if sig_982 = '1' then
				dec_plt2 <= mux_500;
			end if;
			if sig_1132 = '1' then
				dec_plt1 <= mux_498;
			end if;
			if sig_906 = '1' then
				dec_plt <= sig_1289(31 downto 0);
			end if;
			if sig_906 = '1' then
				dec_sl <= sig_1298(31 downto 0);
			end if;
			if sig_897 = '1' then
				dec_rlt <= sig_1298(30 downto 0);
			end if;
			if sig_982 = '1' then
				dec_rlt2 <= mux_490;
			end if;
			if sig_1132 = '1' then
				dec_rlt1 <= mux_488;
			end if;
			if sig_1014 = '1' then
				dec_al2 <= mux_486;
			end if;
			if sig_992 = '1' then
				dec_al1 <= mux_484;
			end if;
			if sig_913 = '1' then
				dl <= sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31) & sig_1281(31 downto 15);
			end if;
			if sig_1014 = '1' then
				dec_nbh <= mux_480;
			end if;
			if sig_897 = '1' then
				dec_dh <= sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 15);
			end if;
			if sig_1030 = '1' then
				dec_nbl <= mux_476;
			end if;
			if sig_1258 = '1' then
				dec_rh2 <= mux_474;
			end if;
			if sig_981 = '1' then
				dec_rh1 <= mux_472;
			end if;
			if sig_1026 = '1' then
				dec_ah2 <= mux_470;
			end if;
			if sig_1058 = '1' then
				dec_ah1 <= mux_468;
			end if;
			if sig_894 = '1' then
				dec_ph <= sig_1298(31 downto 0);
			end if;
			if sig_894 = '1' then
				dec_sh <= sig_1289(31 downto 0);
			end if;
			if sig_1258 = '1' then
				dec_ph2 <= mux_462;
			end if;
			if sig_981 = '1' then
				dec_ph1 <= mux_460;
			end if;
			if sig_975 = '1' then
				abs_m_3 <= mux_458;
			end if;
			if sig_1232 = '1' then
				filtep_pl_14 <= mux_456;
			end if;
			if sig_965 = '1' then
				quantl_el_16 <= el(31);
			end if;
			if sig_867 = '1' then
				quantl_detl_17 <= detl;
			end if;
			if sig_1063 = '1' then
				quantl_ril_18 <= or_669;
			end if;
			if sig_900 = '1' then
				quantl_mil_19 <= mux_448;
			end if;
			if sig_1024 = '1' then
				quantl_wd_20 <= abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3(31) & abs_m_3;
			end if;
			if sig_1158 = '1' then
				quantl_decis_21 <= sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31) & sig_1304(31 downto 15);
			end if;
			if sig_1106 = '1' then
				logscl_nbl_27 <= mux_440;
			end if;
			if sig_1060 = '1' then
				logscl_wd_28 <= mux_438;
			end if;
			if sig_1067 = '1' then
				scalel_wd3_35 <= sig_1295(28 downto 0);
			end if;
			if sig_1259 = '1' then
				uppol2_wd4_42 <= mux_434;
			end if;
			if sig_1165 = '1' then
				uppol2_apl2_43 <= mux_432;
			end if;
			if sig_1259 = '1' then
				uppol1_wd2_51 <= mux_430;
			end if;
			if sig_1028 = '1' then
				uppol1_wd3_52 <= sig_1302(31 downto 0);
			end if;
			if sig_1134 = '1' then
				uppol1_apl1_53 <= mux_426;
			end if;
			if sig_1141 = '1' then
				logsch_nbh_57 <= mux_424;
			end if;
			if sig_1148 = '1' then
				logsch_wd_58 <= mux_422;
			end if;
			if sig_867 = '1' then
				encode_xin1_61 <= sig_1296;
			end if;
			if sig_867 = '1' then
				encode_xin2_62 <= sig_1297;
			end if;
			if sig_1225 = '1' then
				encode_xa_67 <= mux_416;
			end if;
			if sig_1225 = '1' then
				encode_xb_68 <= mux_414;
			end if;
			if sig_1152 = '1' then
				encode_decis_69 <= sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31) & sig_1291(31 downto 12);
			end if;
			if sig_913 = '1' then
				decode_input_98 <= sig_1294(31 downto 2);
			end if;
			if sig_1144 = '1' then
				decode_xa1_100 <= mux_406;
			end if;
			if sig_1144 = '1' then
				decode_xa2_101 <= mux_404;
			end if;
			if sig_1138 = '1' then
				augh_main_i_132 <= mux_372;
			end if;
			if sig_996 = '1' then
				encode_ret0_136 <= or_699 & quantl_ril_18(5 downto 0);
			end if;
			if sig_1258 = '1' then
				dec_del_dhx_reg0 <= mux_338;
			end if;
			if sig_1258 = '1' then
				dec_del_dhx_reg1 <= mux_336;
			end if;
			if sig_980 = '1' then
				dec_del_bph_reg0 <= mux_326;
			end if;
			if sig_979 = '1' then
				dec_del_bph_reg1 <= mux_324;
			end if;
			if sig_977 = '1' then
				dec_del_bph_reg2 <= mux_322;
			end if;
			if sig_1164 = '1' then
				dec_del_bph_reg3 <= mux_320;
			end if;
			if sig_978 = '1' then
				dec_del_bph_reg4 <= mux_318;
			end if;
			if sig_1170 = '1' then
				dec_del_bph_reg5 <= mux_316;
			end if;
			if sig_982 = '1' then
				dec_del_dltx_reg0 <= mux_310;
			end if;
			if sig_982 = '1' then
				dec_del_dltx_reg1 <= mux_308;
			end if;
			if sig_1264 = '1' then
				dec_del_bpl_reg0 <= mux_298;
			end if;
			if sig_1051 = '1' then
				dec_del_bpl_reg1 <= mux_296;
			end if;
			if sig_1267 = '1' then
				dec_del_bpl_reg2 <= mux_294;
			end if;
			if sig_1052 = '1' then
				dec_del_bpl_reg3 <= mux_292;
			end if;
			if sig_1173 = '1' then
				dec_del_bpl_reg4 <= mux_290;
			end if;
			if sig_1050 = '1' then
				dec_del_bpl_reg5 <= mux_288;
			end if;
			if sig_1116 = '1' then
				delay_bph_reg0 <= mux_286;
			end if;
			if sig_1279 = '1' then
				delay_bph_reg1 <= mux_284;
			end if;
			if sig_1111 = '1' then
				delay_bph_reg2 <= mux_282;
			end if;
			if sig_1110 = '1' then
				delay_bph_reg3 <= mux_280;
			end if;
			if sig_1113 = '1' then
				delay_bph_reg4 <= mux_278;
			end if;
			if sig_1114 = '1' then
				delay_bph_reg5 <= mux_276;
			end if;
			if sig_998 = '1' then
				delay_dhx_reg0 <= mux_274;
			end if;
			if sig_998 = '1' then
				delay_dhx_reg1 <= mux_272;
			end if;
			if sig_1151 = '1' then
				delay_dltx_reg0 <= mux_262;
			end if;
			if sig_1151 = '1' then
				delay_dltx_reg1 <= mux_260;
			end if;
			if sig_1131 = '1' then
				delay_bpl_reg0 <= mux_250;
			end if;
			if sig_1128 = '1' then
				delay_bpl_reg1 <= mux_248;
			end if;
			if sig_1126 = '1' then
				delay_bpl_reg2 <= mux_246;
			end if;
			if sig_1124 = '1' then
				delay_bpl_reg3 <= mux_244;
			end if;
			if sig_1127 = '1' then
				delay_bpl_reg4 <= mux_242;
			end if;
			if sig_1130 = '1' then
				delay_bpl_reg5 <= mux_240;
			end if;
			if sig_1006 = '1' then
				accumc_reg0 <= mux_238;
			end if;
			if sig_1006 = '1' then
				accumc_reg1 <= mux_236;
			end if;
			if sig_1006 = '1' then
				accumc_reg2 <= mux_234;
			end if;
			if sig_1006 = '1' then
				accumc_reg3 <= mux_232;
			end if;
			if sig_1006 = '1' then
				accumc_reg4 <= mux_230;
			end if;
			if sig_1006 = '1' then
				accumc_reg5 <= mux_228;
			end if;
			if sig_1006 = '1' then
				accumc_reg6 <= mux_226;
			end if;
			if sig_1006 = '1' then
				accumc_reg7 <= mux_224;
			end if;
			if sig_1006 = '1' then
				accumc_reg8 <= mux_222;
			end if;
			if sig_1006 = '1' then
				accumc_reg9 <= mux_220;
			end if;
			if sig_1006 = '1' then
				accumc_reg10 <= mux_218;
			end if;
			if sig_1006 = '1' then
				accumd_reg0 <= mux_216;
			end if;
			if sig_1006 = '1' then
				accumd_reg1 <= mux_214;
			end if;
			if sig_1006 = '1' then
				accumd_reg2 <= mux_212;
			end if;
			if sig_1006 = '1' then
				accumd_reg3 <= mux_210;
			end if;
			if sig_1006 = '1' then
				accumd_reg4 <= mux_208;
			end if;
			if sig_1006 = '1' then
				accumd_reg5 <= mux_206;
			end if;
			if sig_1006 = '1' then
				accumd_reg6 <= mux_204;
			end if;
			if sig_1006 = '1' then
				accumd_reg7 <= mux_202;
			end if;
			if sig_1006 = '1' then
				accumd_reg8 <= mux_200;
			end if;
			if sig_1006 = '1' then
				accumd_reg9 <= mux_198;
			end if;
			if sig_1006 = '1' then
				accumd_reg10 <= mux_196;
			end if;
			if sig_1176 = '1' then
				tqmf_reg8 <= mux_194;
			end if;
			if sig_1176 = '1' then
				tqmf_reg9 <= mux_192;
			end if;
			if sig_1176 = '1' then
				tqmf_reg10 <= mux_190;
			end if;
			if sig_1176 = '1' then
				tqmf_reg11 <= mux_188;
			end if;
			if sig_1176 = '1' then
				tqmf_reg12 <= mux_186;
			end if;
			if sig_1176 = '1' then
				tqmf_reg13 <= mux_184;
			end if;
			if sig_1176 = '1' then
				tqmf_reg14 <= mux_182;
			end if;
			if sig_1176 = '1' then
				tqmf_reg15 <= mux_180;
			end if;
			if sig_1176 = '1' then
				tqmf_reg16 <= mux_178;
			end if;
			if sig_1176 = '1' then
				tqmf_reg17 <= mux_176;
			end if;
			if sig_1176 = '1' then
				tqmf_reg18 <= mux_174;
			end if;
			if sig_1176 = '1' then
				tqmf_reg19 <= mux_172;
			end if;
			if sig_1176 = '1' then
				tqmf_reg20 <= mux_170;
			end if;
			if sig_1176 = '1' then
				tqmf_reg21 <= mux_168;
			end if;
			if sig_1176 = '1' then
				tqmf_reg22 <= mux_166;
			end if;
			if sig_1176 = '1' then
				tqmf_reg23 <= mux_164;
			end if;
		end if;
	end process;

	-- Remaining signal assignments
	-- Those who are not assigned by component instantiation

	sig_clock <= clock;
	sig_reset <= reset;
	augh_test_23 <= sig_1300;
	augh_test_24 <= sig_1300;
	sig_start <= start;
	augh_test_135 <= sig_1300;
	augh_test_137 <= sig_1300;
	augh_test_138 <= sig_1300;
	sig_1319 <= uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43(31) & uppol2_apl2_43;

	-- Remaining top-level ports assignments
	-- Those who are not assigned by component instantiation

	stdin_rdy <= sig_1221;
	stdout_data <= write32_val_1;

end architecture;
