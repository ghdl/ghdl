entity simple is
end simple;

architecture behav of simple is
begin
  assert false report "Hello";
end behav;
