package badrng is
    signal Sht : bit_vector(2 downtonatural range 0 to 7;
end badrng;
