entity var1 is
end;

use work.pkg.all;

architecture behav of var1 is
begin
  process
   variable v : rec_4;
  begin
   wait;
  end process;
end behav;
