-- comments before design units :ctx1:
--:ctx1: might be multiline
context ctx1 is
end context;
