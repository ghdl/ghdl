library ieee;
use ieee.std_logic_1164.all;

entity underscore1 is
  constant v : std_logic_vector := b"_10";
end;
