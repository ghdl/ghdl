
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc195.vhd,v 1.2 2001-10-26 16:30:14 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s00b00x00p11n01i00195ent IS
END c03s00b00x00p11n01i00195ent;

ARCHITECTURE c03s00b00x00p11n01i00195arch OF c03s00b00x00p11n01i00195ent IS
  type       T1 is array (0 to 31) of BIT;
  subtype    T2 is integer range 2 to 20;
  signal    S1 : T2 ;
BEGIN
  TESTING: PROCESS
  BEGIN
    S1 <= 25 after 10 ns; 
    wait for 20 ns;
    assert NOT(S1 = 25)
      report "***PASSED TEST: c03s00b00x00p11n01i00195"
      severity NOTE;
    assert ( S1 = 25 )
      report "***FAILED TEST: c03s00b00x00p11n01i00195 - Value doesn't belong to the range of the subtype of the object." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s00b00x00p11n01i00195arch;
