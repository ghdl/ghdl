library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package TestPkg is

end package TestPkg ; 
