entity r is
end;
