package--
function(0is
while()0X';