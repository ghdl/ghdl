-- Author:  Patrick Lehmann
-- License: MIT
--
-- undocumented
--
context StopWatch_ctx is
	library lib_Utilities;
	context lib_Utilities.Utilities_pkg;

	use work.StopWatch_pkg.all;
end context;
