package p is
  --  Comment for :rec:
  type rec is record
    a : bit;
    b : bit;
  end record;
end p;
