
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1804.vhd,v 1.2 2001-10-26 16:29:43 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c07s01b00x00p06n01i01804ent IS
END c07s01b00x00p06n01i01804ent;

ARCHITECTURE c07s01b00x00p06n01i01804arch OF c07s01b00x00p06n01i01804ent IS

BEGIN
  TESTING: PROCESS
    variable x : integer := 0;
    variable y : integer := 2;
    variable z : integer := 5;
  BEGIN
    x := y * 10 * z;  -- No_failure_here
    assert NOT( x=100 )
      report "***PASSED TEST: c07s01b00x00p06n01i01804"
      severity NOTE;
    assert ( x=100 )
      report "***FAILED TEST: c07s01b00x00p06n01i01804 - The term must be factor or a sequence of factors combined with multiplying operators."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c07s01b00x00p06n01i01804arch;
