
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1138.vhd,v 1.2 2001-10-26 16:29:39 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c06s05b00x00p05n02i01138ent IS
END c06s05b00x00p05n02i01138ent;

ARCHITECTURE c06s05b00x00p05n02i01138arch OF c06s05b00x00p05n02i01138ent IS
  signal T1 : boolean;
BEGIN
  TESTING: PROCESS
    variable B : Bit_vector (1 to 10) := B"01010_10101";
  BEGIN
    if B(1 to 2) = B"01"  then
      T1 <= TRUE;
    else
      T1 <= FALSE;
    end if;
    wait for 1 ns;
    assert NOT(T1=TRUE)
      report "***PASSED TEST: c06s05b00x00p05n02i01138"
      severity NOTE;
    assert (T1=TRUE)
      report "***FAILED TEST: c06s05b00x00p05n02i01138 - The prefix and the discrete range of the slice is not correctly evaluated."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c06s05b00x00p05n02i01138arch;
