package data_pkg is
  type word_vector is array (natural range <>) of
      Natural;

  constant data : word_vector := (
    16#56f8f7d0#, 16#6dee3844#, 16#6ed60624#, 16#617fd1e0#, 
    16#20053fe6#, 16#200b3301#, 16#74a469d5#, 16#2791b468#, 
    16#2a36168d#, 16#3d06b618#, 16#3531c529#, 16#59b86d4b#, 
    16#38392b2d#, 16#0048d40c#, 16#015447e5#, 16#048382d3#, 
    16#19ca235a#, 16#44b8edec#, 16#75c052d6#, 16#7339660a#, 
    16#4a47b6ce#, 16#3f3af14c#, 16#4d5dd733#, 16#48bd0b2d#, 
    16#49497750#, 16#5415889a#, 16#5ad38e67#, 16#74e47c34#, 
    16#5e974b6e#, 16#6b3026d2#, 16#41fd020e#, 16#5135fdb3#, 
    16#0db780ba#, 16#614d9c7e#, 16#18c1d4c0#, 16#3de1e866#, 
    16#3987cc45#, 16#182937b3#, 16#0510fa65#, 16#7361a5ce#, 
    16#19e2df54#, 16#72356dc7#, 16#232e0a67#, 16#53741bfa#, 
    16#36456b90#, 16#4e626d08#, 16#3970562a#, 16#58fb0379#, 
    16#411eabee#, 16#0261ba7b#, 16#4e07878a#, 16#33458e41#, 
    16#3b82ca1a#, 16#4ccfc0e9#, 16#356b5f7e#, 16#3051d779#, 
    16#338ad77b#, 16#460ca8b7#, 16#66724dfe#, 16#24333e95#, 
    16#5530f83d#, 16#4b70cf86#, 16#6efeda26#, 16#62cd22ea#, 
    16#4f15a22a#, 16#49725a8f#, 16#3c6b4d80#, 16#73897db0#, 
    16#7ee49383#, 16#5f15708e#, 16#53159cba#, 16#21667155#, 
    16#1117d4dd#, 16#3b55f182#, 16#50de52ef#, 16#1ea017d3#, 
    16#6e2d90b2#, 16#6190f475#, 16#76baa3ce#, 16#2391e255#, 
    16#69919317#, 16#5e738aa3#, 16#5d71ec39#, 16#3f55d989#, 
    16#056dc86f#, 16#0ed98f1f#, 16#793a13fc#, 16#51a3106c#, 
    16#18aa7637#, 16#602529b8#, 16#4d81440c#, 16#7204dc43#, 
    16#53990a6d#, 16#65745255#, 16#176f333a#, 16#5603e66a#, 
    16#391d0c3d#, 16#00071cc4#, 16#64d51d48#, 16#796ad40b#, 
    16#445b6e3d#, 16#0f0a8ed6#, 16#38fffd86#, 16#17c1316b#, 
    16#1bf1ebfb#, 16#2e1d88ff#, 16#47bee4ee#, 16#4e8b6fde#, 
    16#62c739ed#, 16#5aca0d1e#, 16#2530ffe3#, 16#4d51b90c#, 
    16#795a86a5#, 16#3e354605#, 16#24268c5e#, 16#6ec8993b#, 
    16#432d1f9a#, 16#33606edf#, 16#2ad49328#, 16#5da953e9#, 
    16#4fdbf363#, 16#2b191322#, 16#7d560358#, 16#5aad74cb#, 
    16#2314d477#, 16#67d73ddf#, 16#053b6780#, 16#68a071dc#, 
    16#0b6bbd91#, 16#5d3eaa7d#, 16#5344f982#, 16#7767d15c#, 
    16#57f7ad77#, 16#68d5ad0f#, 16#5018defb#, 16#7be3b5de#, 
    16#39ca0f9f#, 16#141103f8#, 16#4fee454c#, 16#48dbbef2#, 
    16#16349958#, 16#271d5150#, 16#71399dfe#, 16#5c42c326#, 
    16#7675f543#, 16#5165199b#, 16#7b731780#, 16#23e0e260#, 
    16#17afa847#, 16#5acd3e24#, 16#4daaf2b3#, 16#13152b35#, 
    16#122ea92b#, 16#1e8eba51#, 16#5fb92e55#, 16#56a8fec4#, 
    16#5634e05e#, 16#143c5ba4#, 16#1e6cfc95#, 16#68f7cbe5#, 
    16#76a95004#, 16#6913c731#, 16#5d2ba93c#, 16#35672599#, 
    16#688c41f6#, 16#02c93bfb#, 16#2fbeae2e#, 16#7032098d#, 
    16#2a414101#, 16#165efcd3#, 16#68f5f326#, 16#3b257de1#, 
    16#6a8c0a66#, 16#08ed5bcd#, 16#208ca8bd#, 16#27066e49#, 
    16#0c7c5bc0#, 16#30582d3a#, 16#79080117#, 16#08cc54a3#, 
    16#1c45e61e#, 16#080ee934#, 16#548a34fd#, 16#2ac69d96#, 
    16#136e5d8a#, 16#15997b07#, 16#1bc8cf68#, 16#36ac8711#, 
    16#1999377b#, 16#49db3e29#, 16#1c0b53e0#, 16#50b67a45#, 
    16#7f0db46f#, 16#74f89f26#, 16#286e2529#, 16#46574069#, 
    16#36aaf8ac#, 16#40966e86#, 16#5bbb7b4d#, 16#60da14a6#, 
    16#6a381ac7#, 16#2caf4c9d#, 16#36f4ae85#, 16#2063fd2e#, 
    16#1bdbe983#, 16#5c8fccd6#, 16#1988bd45#, 16#79d6201e#, 
    16#21636cda#, 16#3b7be5f0#, 16#1bb4fa48#, 16#121d2bf8#, 
    16#4cd3d6e5#, 16#2857a4db#, 16#27b9ab01#, 16#6bf797fe#, 
    16#49a65211#, 16#0d44b24a#, 16#7edf9a73#, 16#1676fb2d#, 
    16#32321909#, 16#23cc9149#, 16#37e5a46f#, 16#1da6ba5f#, 
    16#37872a46#, 16#2cb92014#, 16#0442a250#, 16#620042d6#, 
    16#116e428d#, 16#3e9f53cc#, 16#5a4a43a6#, 16#2290c175#, 
    16#7578c1ae#, 16#5db958e3#, 16#466b202c#, 16#2b718592#, 
    16#3b4f1367#, 16#18567871#, 16#1f212009#, 16#20b1bb1f#, 
    16#4967535e#, 16#4177ee95#, 16#47bdff3c#, 16#450c44d8#, 
    16#47ac748d#, 16#384a5d38#, 16#109d53ce#, 16#3b5e594f#, 
    16#3b261875#, 16#50131c16#, 16#29bfce20#, 16#22a1cb8d#, 
    16#788c5553#, 16#7befe74b#, 16#1a1abff1#, 16#458ecb93#, 
    16#2e0bb25c#, 16#0f33c86c#, 16#21d2215d#, 16#67d8bd0d#, 
    16#29d2d6c8#, 16#2a0642d9#, 16#64e51b00#, 16#72aa9215#, 
    16#7b6003ff#, 16#3003674a#, 16#61f5542e#, 16#66dce744#, 
    16#1e6afce1#, 16#191329b8#, 16#3def1315#, 16#7cd937b9#, 
    16#76c3b12e#, 16#5acee9d9#, 16#22f0071e#, 16#06c8ec01#, 
    16#0e8cefd5#, 16#421d3c32#, 16#57f28e9f#, 16#45e03422#, 
    16#241d1772#, 16#55c6e83d#, 16#1e3b9f41#, 16#56ceb1ee#, 
    16#24b50b14#, 16#120bc455#, 16#66fdea7c#, 16#3e6080a1#, 
    16#19053cad#, 16#1987fc79#, 16#713bceed#, 16#56d3dcfe#, 
    16#14beb12b#, 16#348ebd1d#, 16#77bde7f0#, 16#0adbb01e#, 
    16#0071d432#, 16#2985797f#, 16#1d20c29d#, 16#1a4af25e#, 
    16#5146cdbc#, 16#07eed480#, 16#4edcccb7#, 16#270762a9#, 
    16#7678f3db#, 16#6b45454b#, 16#1b93046f#, 16#2ef023f7#, 
    16#55e8dbfa#, 16#7f8cb85f#, 16#628fa6b3#, 16#05efb9dd#, 
    16#3de62c05#, 16#0f6a4fe8#, 16#34d15a7e#, 16#42b4c25b#, 
    16#33c084bf#, 16#062fc9b0#, 16#1b6bdf55#, 16#405c63e0#, 
    16#5157bb23#, 16#414f84d2#, 16#4f78eb50#, 16#375be80e#, 
    16#5e3b08d9#, 16#291d0e2f#, 16#7dcacf1d#, 16#1dc3a484#, 
    16#2304693b#, 16#03187825#, 16#30cacce6#, 16#7c987679#, 
    16#49b45cc8#, 16#4b0b4461#, 16#2c6f7b87#, 16#1e982ad0#, 
    16#789cf214#, 16#2566768c#, 16#72e6a3da#, 16#1f0262d3#, 
    16#194b5b06#, 16#2b19cbfb#, 16#772b2c8d#, 16#3540ffef#, 
    16#2b003d97#, 16#0419aa23#, 16#79c325da#, 16#2775313b#, 
    16#0f0692eb#, 16#0073e0a0#, 16#0290aeef#, 16#15e2078c#, 
    16#22480767#, 16#41520845#, 16#1a13f538#, 16#33954b20#, 
    16#78dcae8e#, 16#448c3836#, 16#1e4451fb#, 16#364cabb9#, 
    16#2f42d973#, 16#1cf46314#, 16#2f13afed#, 16#4c6cd961#, 
    16#799e4a12#, 16#156dfc1b#, 16#6b8aa648#, 16#6f8975e0#, 
    16#21a9c8b7#, 16#5c8bf777#, 16#59c8d814#, 16#70490f68#, 
    16#03add532#, 16#2bb1e36f#, 16#0b0bb981#, 16#5c2e0d17#, 
    16#2b4db850#, 16#0ce24274#, 16#5ed2aa3d#, 16#6b671a14#, 
    16#03027153#, 16#7854842d#, 16#0a01b4fc#, 16#6191da20#, 
    16#44d43b36#, 16#55584f90#, 16#364ea359#, 16#1d7a2f3a#, 
    16#5b3ce52e#, 16#5c102f8d#, 16#7516d7ee#, 16#455d447f#, 
    16#3784a1d9#, 16#2780c979#, 16#220e0cbe#, 16#07b30842#, 
    16#10caa080#, 16#5511a525#, 16#55833137#, 16#1c239b35#, 
    16#24901caa#, 16#01fae8e6#, 16#7a86c13e#, 16#3e334c49#, 
    16#0acf5b14#, 16#62e61cf1#, 16#6c804b72#, 16#2923dad6#, 
    16#52667409#, 16#1023e592#, 16#77eeca14#, 16#284d1480#, 
    16#43a71018#, 16#5db67e47#, 16#47a4513a#, 16#6e863287#, 
    16#1a3da2e9#, 16#0f7a43e4#, 16#452cefe4#, 16#719c7987#, 
    16#73923963#, 16#3a83b1c9#, 16#35d28e02#, 16#30e65a89#, 
    16#1b29499e#, 16#02e0b650#, 16#3ed4df9d#, 16#31315d7e#, 
    16#1228a1fa#, 16#6d06f9f1#, 16#76aaa090#, 16#7812c415#, 
    16#29dd1228#, 16#08b344b3#, 16#35dae9a7#, 16#50343668#, 
    16#2fd7bca0#, 16#54a8aa33#, 16#29b46756#, 16#629914ff#, 
    16#230ca0aa#, 16#717c424b#, 16#79e10ae2#, 16#57207af3#, 
    16#13b36a87#, 16#78c71cb0#, 16#747e0480#, 16#336480a5#, 
    16#68cee5e0#, 16#467b0ffb#, 16#1e2c844b#, 16#5c4dc53f#, 
    16#50f20c8a#, 16#69f49c29#, 16#08af735c#, 16#7552eaa9#, 
    16#34fff369#, 16#0bc34cfb#, 16#3463b947#, 16#5691ba41#, 
    16#337f9288#, 16#062e015a#, 16#37440a0d#, 16#7c92ded2#, 
    16#421ca91f#, 16#50b6eb2d#, 16#4e9b5f1e#, 16#4ac1cbc6#, 
    16#64d6fd0d#, 16#7638df8c#, 16#7b3d6bf7#, 16#6375d6d5#, 
    16#275a7802#, 16#2d8f115c#, 16#09fe3b88#, 16#2c54b7de#, 
    16#0ea40779#, 16#4e795a57#, 16#06ca0179#, 16#6c6122ae#, 
    16#78f69fdd#, 16#6d250285#, 16#2be6759d#, 16#12809ba6#, 
    16#031e2012#, 16#4cc034b5#, 16#4af54907#, 16#76d60004#, 
    16#47e7934c#, 16#684bc376#, 16#1cba80ec#, 16#4c6dcbfc#, 
    16#407bd0a9#, 16#0cb74076#, 16#3aa53ba2#, 16#26a2d7c3#, 
    16#0b6b41ac#, 16#411cacc1#, 16#0d661f7d#, 16#79e45873#, 
    16#009bfd85#, 16#24fd3f46#, 16#04e25e0d#, 16#786a280c#, 
    16#14c8e7b0#, 16#339e4280#, 16#02971b52#, 16#4bfbf050#, 
    16#2634c43a#, 16#3a8226ab#, 16#42fa55b8#, 16#2971d073#, 
    16#6b5f0441#
    );
end data_pkg;
