library ieee;
use ieee.std_logic_1164.all;

package repro is
  alias reg_Acc is "0111";
end repro;
