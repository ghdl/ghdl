package function(0is if X�X';