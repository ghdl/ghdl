package function return g.b of