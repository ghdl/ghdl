
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc848.vhd,v 1.2 2001-10-26 16:30:28 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c01s03b01x00p09n01i00848ent IS
  port ( PT : Boolean );
END c01s03b01x00p09n01i00848ent;

ARCHITECTURE c01s03b01x00p09n01i00848arch OF c01s03b01x00p09n01i00848ent IS

BEGIN

  BD : block
    component comp1
    end component ;
  begin
    CIS : comp1;
    BD_nested : block
    begin
      process
      begin
        null;
        wait;
      End process;
    end block;
  end block BD ;

  TESTING: PROCESS
  BEGIN
    assert FALSE 
      report "***FAILED TEST: c01s03b01x00p09n01i00848 - Invalid block specification."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c01s03b01x00p09n01i00848arch;

configuration c01s03b01x00p09n01i00848cfg of c01s03b01x00p09n01i00848ent is
  for c01s03b01x00p09n01i00848arch
    for CIS  -- Failure_here
      -- ERROR: the CIS is not a declared block in the declarative region.
    end for ;
    for BD_nested  -- failure_here
      -- ERROR :: BD_nested is not a block label in the related declarative region.
    end for;
  end for;
end c01s03b01x00p09n01i00848cfg;
