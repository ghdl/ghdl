package p is
  type rec is record
    a : bit;
    --  Comment for the first element :b:
    b : bit;
  end record;
end p;
