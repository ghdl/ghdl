library IEEE;
use IEEE.std_logic_1164.all;

package protocol_pkg is
    type T_ARRAY is array (NATURAL range <>) of STD_LOGIC_VECTOR;
end protocol_pkg;
