entity e is
  generic(type t);
  signal w:integer range 0 to t;
end;
