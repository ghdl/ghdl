
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc100.vhd,v 1.2 2001-10-26 16:29:38 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

package c04s03b02x00p29n06i00100pkg is
  type int_1 is range 1 to 32;
  attribute pin_number : int_1;
end c04s03b02x00p29n06i00100pkg;

use work.c04s03b02x00p29n06i00100pkg.all;
ENTITY c04s03b02x00p29n06i00100ent IS
  port ( P2 : out bit) ;
  attribute pin_number of P2 : signal is 1;
END c04s03b02x00p29n06i00100ent;

ARCHITECTURE c04s03b02x00p29n06i00100arch OF c04s03b02x00p29n06i00100ent IS

BEGIN
  TESTING: PROCESS
    variable pn : int_1;
  BEGIN
    pn := 1;
    assert NOT( P2'pin_number = pn )
      report "***PASSED TEST: c04s03b02x00p29n06i00100"      severity NOTE;
    assert ( P2'pin_number = pn )
      report "***FAILED TEST: c04s03b02x00p29n06i00100 - Reading user defined attributes of interface elements of mode 'out' should be permitted."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c04s03b02x00p29n06i00100arch;
