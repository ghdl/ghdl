
-- Copyright (C) 2002 Morgan Kaufmann Publishers, Inc

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

entity inline_10a is

end entity inline_10a;


----------------------------------------------------------------


architecture test of inline_10a is

  -- code from book:

  type stick_position is (down, center, up);

  -- end of code from book

  signal throttle : stick_position;

begin


  process_3_a : process (throttle) is

    variable speed : integer := 0;
    constant decrement : integer := 1;
    constant increment : integer := 1;

  begin

    -- code from book:

    case throttle is
      when down =>
        speed := speed - decrement;
      when up =>
        speed := speed + increment;
      when center =>
        null; -- no change to speed
    end case;

    -- end of code from book

  end process process_3_a;


  stimulus : process is
  begin
    throttle <= down after 10 ns, center after 20 ns, up after 30 ns;
    wait;
  end process stimulus;


end architecture test;
