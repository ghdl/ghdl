package p2 is
  -- comments in design units (python doc-string style) :fail:

  constant c : natural := 5;
end package;
