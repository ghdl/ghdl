
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1909.vhd,v 1.2 2001-10-26 16:29:43 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c07s02b00x00p09n03i01909ent IS
END c07s02b00x00p09n03i01909ent;

ARCHITECTURE c07s02b00x00p09n03i01909arch OF c07s02b00x00p09n03i01909ent IS
  signal Q     : BIT := '1';
  signal R     : BIT := '0';
  signal S     : BIT := '1';
  signal PP,P2 : BIT := '1' ;
  signal R1    : BIT;
BEGIN
  TESTING: PROCESS
  BEGIN
    R1 <= ((Q and S) or R) and (P2 and PP) ;
    wait for 5 ns;
    assert NOT( R1 = '1' )
      report "***PASSED TEST: c07s02b00x00p09n03i01909"
      severity NOTE;
    assert ( R1 = '1' )
      report "***FAILED TEST: c07s02b00x00p09n03i01909 - The parentheses can be used to control the association of operators and operands."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c07s02b00x00p09n03i01909arch;
