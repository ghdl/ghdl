package issue_pkg is

  type t_one_two is (one, two);

end package issue_pkg;
