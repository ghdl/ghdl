
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1547.vhd,v 1.2 2001-10-26 16:29:42 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c08s09b00x00p10n01i01547ent IS
END c08s09b00x00p10n01i01547ent;

ARCHITECTURE c08s09b00x00p10n01i01547arch OF c08s09b00x00p10n01i01547ent IS

BEGIN
  TESTING: PROCESS
    type     t_enum1 is (en1, en2, en3, en4) ;
    subtype  st_enum1 is t_enum1 range en4 downto en1 ;
    variable counter : integer := 0;
  BEGIN
    for i in st_enum1 loop
      counter := counter + 1;
    end loop;
    assert NOT(counter=st_enum1'Pos(st_enum1'High)-st_enum1'Pos(st_enum1'Low)+1) 
      report "***PASSED TEST: c08s09b00x00p10n01i01547" 
      severity NOTE;
    assert (counter=st_enum1'Pos(st_enum1'High)-st_enum1'Pos(st_enum1'Low)+1) 
      report "***FAILED TEST: c08s09b00x00p10n01i01547 - The loop is executed once for each of the values in the range." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c08s09b00x00p10n01i01547arch;
