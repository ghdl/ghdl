entity test is
end test;

architecture only of test is
begin  -- only
  doit: process
  begin  -- process
    assert( character'pos(NUL) = 0 ) report "TEST FAILED" severity failure;
    assert ( character'pos(SOH) = 1)  report "TEST FAILED" severity failure;
    assert ( character'pos(STX) = 2)  report "TEST FAILED" severity failure;
    assert ( character'pos(ETX) = 3)  report "TEST FAILED" severity failure;
    assert ( character'pos(EOT) = 4)  report "TEST FAILED" severity failure;
    assert ( character'pos(ENQ) = 5)  report "TEST FAILED" severity failure;
    assert ( character'pos(ACK) = 6)  report "TEST FAILED" severity failure;
    assert ( character'pos(BEL) = 7)  report "TEST FAILED" severity failure;
    assert ( character'pos(BS ) = 8)  report "TEST FAILED" severity failure;
    assert ( character'pos(HT ) = 9)  report "TEST FAILED" severity failure;
    assert ( character'pos(LF ) = 10)  report "TEST FAILED" severity failure;
    assert ( character'pos(VT ) = 11)  report "TEST FAILED" severity failure;
    assert ( character'pos(FF ) = 12)  report "TEST FAILED" severity failure;
    assert ( character'pos(CR ) = 13)  report "TEST FAILED" severity failure;
    assert ( character'pos(SO ) = 14)  report "TEST FAILED" severity failure;
    assert ( character'pos(SI ) = 15)  report "TEST FAILED" severity failure;
    assert ( character'pos(DLE) = 16)  report "TEST FAILED" severity failure;
    assert ( character'pos(DC1) = 17)  report "TEST FAILED" severity failure;
    assert ( character'pos(DC2) = 18)  report "TEST FAILED" severity failure;
    assert ( character'pos(DC3) = 19)  report "TEST FAILED" severity failure;
    assert ( character'pos(DC4) = 20)  report "TEST FAILED" severity failure;
    assert ( character'pos(NAK) = 21)  report "TEST FAILED" severity failure;
    assert ( character'pos(SYN) = 22)  report "TEST FAILED" severity failure;
    assert ( character'pos(ETB) = 23)  report "TEST FAILED" severity failure;
    assert ( character'pos(CAN) = 24)  report "TEST FAILED" severity failure;
    assert ( character'pos(EM ) = 25)  report "TEST FAILED" severity failure;
    assert ( character'pos(SUB) = 26)  report "TEST FAILED" severity failure;
    assert ( character'pos(ESC) = 27)  report "TEST FAILED" severity failure;
    assert ( character'pos(FSP) = 28)  report "TEST FAILED" severity failure;
    assert ( character'pos(GSP) = 29)  report "TEST FAILED" severity failure;
    assert ( character'pos(RSP) = 30)  report "TEST FAILED" severity failure;
    assert ( character'pos(USP) = 31)  report "TEST FAILED" severity failure;
    assert ( character'pos(' ') = 32)  report "TEST FAILED" severity failure;
    assert ( character'pos('!') = 33)  report "TEST FAILED" severity failure;
    assert ( character'pos('"') = 34)  report "TEST FAILED" severity failure;
    assert ( character'pos('#') = 35)  report "TEST FAILED" severity failure;
    assert ( character'pos('$') = 36)  report "TEST FAILED" severity failure;
    assert ( character'pos('%') = 37)  report "TEST FAILED" severity failure;
    assert ( character'pos('&') = 38)  report "TEST FAILED" severity failure;
    assert ( character'pos(''') = 39)  report "TEST FAILED" severity failure;
    assert ( character'pos('(') = 40)  report "TEST FAILED" severity failure;
    assert ( character'pos(')') = 41)  report "TEST FAILED" severity failure;
    assert ( character'pos('*') = 42)  report "TEST FAILED" severity failure;
    assert ( character'pos('+') = 43)  report "TEST FAILED" severity failure;
    assert ( character'pos(',') = 44)  report "TEST FAILED" severity failure;
    assert ( character'pos('-') = 45)  report "TEST FAILED" severity failure;
    assert ( character'pos('.') = 46)  report "TEST FAILED" severity failure;
    assert ( character'pos('/') = 47)  report "TEST FAILED" severity failure;
    assert ( character'pos('0') = 48)  report "TEST FAILED" severity failure;
    assert ( character'pos('1') = 49)  report "TEST FAILED" severity failure;
    assert ( character'pos('2') = 50)  report "TEST FAILED" severity failure;
    assert ( character'pos('3') = 51)  report "TEST FAILED" severity failure;
    assert ( character'pos('4') = 52)  report "TEST FAILED" severity failure;
    assert ( character'pos('5') = 53)  report "TEST FAILED" severity failure;
    assert ( character'pos('6') = 54)  report "TEST FAILED" severity failure;
    assert ( character'pos('7') = 55)  report "TEST FAILED" severity failure;
    assert ( character'pos('8') = 56)  report "TEST FAILED" severity failure;
    assert ( character'pos('9') = 57)  report "TEST FAILED" severity failure;
    assert ( character'pos(':') = 58)  report "TEST FAILED" severity failure;
    assert ( character'pos(';') = 59)  report "TEST FAILED" severity failure;
    assert ( character'pos('<') = 60)  report "TEST FAILED" severity failure;
    assert ( character'pos('=') = 61)  report "TEST FAILED" severity failure;
    assert ( character'pos('>') = 62)  report "TEST FAILED" severity failure;
    assert ( character'pos('?') = 63)  report "TEST FAILED" severity failure;
    assert ( character'pos('@') = 64)  report "TEST FAILED" severity failure;
    assert ( character'pos('A') = 65)  report "TEST FAILED" severity failure;
    assert ( character'pos('B') = 66)  report "TEST FAILED" severity failure;
    assert ( character'pos('C') = 67)  report "TEST FAILED" severity failure;
    assert ( character'pos('D') = 68)  report "TEST FAILED" severity failure;
    assert ( character'pos('E') = 69)  report "TEST FAILED" severity failure;
    assert ( character'pos('F') = 70)  report "TEST FAILED" severity failure;
    assert ( character'pos('G') = 71)  report "TEST FAILED" severity failure;
    assert ( character'pos('H') = 72)  report "TEST FAILED" severity failure;
    assert ( character'pos('I') = 73)  report "TEST FAILED" severity failure;
    assert ( character'pos('J') = 74)  report "TEST FAILED" severity failure;
    assert ( character'pos('K') = 75)  report "TEST FAILED" severity failure;
    assert ( character'pos('L') = 76)  report "TEST FAILED" severity failure;
    assert ( character'pos('M') = 77)  report "TEST FAILED" severity failure;
    assert ( character'pos('N') = 78)  report "TEST FAILED" severity failure;
    assert ( character'pos('O') = 79)  report "TEST FAILED" severity failure;
    assert ( character'pos('P') = 80)  report "TEST FAILED" severity failure;
    assert ( character'pos('Q') = 81)  report "TEST FAILED" severity failure;
    assert ( character'pos('R') = 82)  report "TEST FAILED" severity failure;
    assert ( character'pos('S') = 83)  report "TEST FAILED" severity failure;
    assert ( character'pos('T') = 84)  report "TEST FAILED" severity failure;
    assert ( character'pos('U') = 85)  report "TEST FAILED" severity failure;
    assert ( character'pos('V') = 86)  report "TEST FAILED" severity failure;
    assert ( character'pos('W') = 87)  report "TEST FAILED" severity failure;
    assert ( character'pos('X') = 88)  report "TEST FAILED" severity failure;
    assert ( character'pos('Y') = 89)  report "TEST FAILED" severity failure;
    assert ( character'pos('Z') = 90)  report "TEST FAILED" severity failure;
    assert ( character'pos('[') = 91)  report "TEST FAILED" severity failure;
    assert ( character'pos('\') = 92)  report "TEST FAILED" severity failure;
    assert ( character'pos(']') = 93)  report "TEST FAILED" severity failure;
    assert ( character'pos('^') = 94)  report "TEST FAILED" severity failure;
    assert ( character'pos('_') = 95)  report "TEST FAILED" severity failure;
    assert ( character'pos('`') = 96)  report "TEST FAILED" severity failure;
    assert ( character'pos('a') = 97)  report "TEST FAILED" severity failure;
    assert ( character'pos('b') = 98)  report "TEST FAILED" severity failure;
    assert ( character'pos('c') = 99)  report "TEST FAILED" severity failure;
    assert ( character'pos('d') = 100)  report "TEST FAILED" severity failure;
    assert ( character'pos('e') = 101)  report "TEST FAILED" severity failure;
    assert ( character'pos('f') = 102)  report "TEST FAILED" severity failure;
    assert ( character'pos('g') = 103)  report "TEST FAILED" severity failure;
    assert ( character'pos('h') = 104)  report "TEST FAILED" severity failure;
    assert ( character'pos('i') = 105)  report "TEST FAILED" severity failure;
    assert ( character'pos('j') = 106)  report "TEST FAILED" severity failure;
    assert ( character'pos('k') = 107)  report "TEST FAILED" severity failure;
    assert ( character'pos('l') = 108)  report "TEST FAILED" severity failure;
    assert ( character'pos('m') = 109)  report "TEST FAILED" severity failure;
    assert ( character'pos('n') = 110)  report "TEST FAILED" severity failure;
    assert ( character'pos('o') = 111)  report "TEST FAILED" severity failure;
    assert ( character'pos('p') = 112)  report "TEST FAILED" severity failure;
    assert ( character'pos('q') = 113)  report "TEST FAILED" severity failure;
    assert ( character'pos('r') = 114)  report "TEST FAILED" severity failure;
    assert ( character'pos('s') = 115)  report "TEST FAILED" severity failure;
    assert ( character'pos('t') = 116)  report "TEST FAILED" severity failure;
    assert ( character'pos('u') = 117)  report "TEST FAILED" severity failure;
    assert ( character'pos('v') = 118)  report "TEST FAILED" severity failure;
    assert ( character'pos('w') = 119)  report "TEST FAILED" severity failure;
    assert ( character'pos('x') = 120)  report "TEST FAILED" severity failure;
    assert ( character'pos('y') = 121)  report "TEST FAILED" severity failure;
    assert ( character'pos('z') = 122)  report "TEST FAILED" severity failure;
    assert ( character'pos('{') = 123)  report "TEST FAILED" severity failure;
    assert ( character'pos('|') = 124)  report "TEST FAILED" severity failure;
    assert ( character'pos('}') = 125)  report "TEST FAILED" severity failure;
    assert ( character'pos('~') = 126)  report "TEST FAILED" severity failure;
    assert ( character'pos(DEL) = 127)  report "TEST FAILED" severity failure;
    assert ( character'pos(character'right) = 255)  report "TEST FAILED" severity failure;
    assert (bit'pos('0') = 0)  report "TEST FAILED" severity failure;
    assert (bit'pos('1') = 1)  report "TEST FAILED" severity failure;
    assert (bit'pos(bit'right) = 1)  report "TEST FAILED" severity failure;
    assert (boolean'pos(false) = 0)  report "TEST FAILED" severity failure;
    assert (boolean'pos(true)  = 1)  report "TEST FAILED" severity failure;
    assert (boolean'pos(boolean'right) = 1)  report "TEST FAILED" severity failure;
    assert (severity_level'pos(NOTE)    = 0)  report "TEST FAILED" severity failure;
    assert (severity_level'pos(WARNING) = 1)  report "TEST FAILED" severity failure;
    assert (severity_level'pos(ERROR)   = 2)  report "TEST FAILED" severity failure;
    assert (severity_level'pos(FAILURE) = 3)  report "TEST FAILED" severity failure;
    assert ( severity_level'pos(severity_level'right) = 3 ) report "TEST FAILED" severity failure;
    report "TEST PASSED";
    wait;
  end process;
end only;
