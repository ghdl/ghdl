
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc271.vhd,v 1.2 2001-10-26 16:30:21 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s01b03x00p06n01i00271ent IS
END c03s01b03x00p06n01i00271ent;

ARCHITECTURE c03s01b03x00p06n01i00271arch OF c03s01b03x00p06n01i00271ent IS
  type GLORIA is range 1 to 6
    units
      PRIM;
      SEC1 = 6 PRIM;
      SEC2 = 36 SEC1;  -- Failure_here
      -- ERROR - SEMANTICS ERROR: Position Number of sec2 exceeds
      -- range of physical type
    end units;
BEGIN
  TESTING: PROCESS
    variable temp : GLORIA := 10 PRIM;
  BEGIN
    assert FALSE 
      report "***FAILED TEST: c03s01b03x00p06n01i00271 - Position number exceeds range of physical type."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s01b03x00p06n01i00271arch;
