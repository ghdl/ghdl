
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc3182.vhd,v 1.2 2001-10-26 16:29:52 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c14s01b00x00p116n01i03182ent IS
END c14s01b00x00p116n01i03182ent;

ARCHITECTURE c14s01b00x00p116n01i03182arch OF c14s01b00x00p116n01i03182ent IS

  constant C : INTEGER := 1;
--
  type t2 is array(c to c + c, 1 to 10) of integer;
  
-- transitive cases
  type t3 is array(t2'range(1), t2'reverse_range(2)) of integer;
  
-- 'Range (of two-dimensional array type)
  type rt311 is range t3'range(1);
  type rt312 is range t3'range(2);

BEGIN
  TESTING: PROCESS
  BEGIN
    wait for 10 ns;
    assert NOT(    rt311'LEFT = rt311(c)   and
                   rt311'RIGHT= rt311(c+c)   and
                   rt312'LEFT = rt312(10)   and
                   rt312'RIGHT= rt312(1)   )
      report "***PASSED TEST: c14s01b00x00p116n01i03182"
      severity NOTE;
    assert (    rt311'LEFT = rt311(c)   and
                rt311'RIGHT= rt311(c+c)   and
                rt312'LEFT = rt312(10)   and
                rt312'RIGHT= rt312(1)   )
      report "***FAILED TEST: c14s01b00x00p116n01i03182 - Predefined attribute range test failed."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c14s01b00x00p116n01i03182arch;
