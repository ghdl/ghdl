architecture@for(""x""4000000000x"