
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2541.vhd,v 1.2 2001-10-26 16:30:19 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c07s03b05x00p14n01i02541ent IS
END c07s03b05x00p14n01i02541ent;

ARCHITECTURE c07s03b05x00p14n01i02541arch OF c07s03b05x00p14n01i02541ent IS

BEGIN
  TESTING: PROCESS
    type X1 is  range 1.0 to 100.0 ;
    type X2 is  range 1.0 to 100.0 ;
    type I1 is  range 1   to 1000000;
    type I2 is  range 1   to 10000000 ;
    variable RE1 : X1 ;
    variable RE2 : X2 ;
    variable IN1 : I1 ;
    variable IN2 : I2 ;
  BEGIN
    RE2 := RE2 * RE1 ;  -- Failure_here
    -- ERROR: TYPE CONVERSION CANNOT OCCUR ON AN OPERAND OF ANY TYPE BUT
    -- UNIVERSAL INTEGER OR UNIVERSAL REAL.
    assert FALSE 
      report "***FAILED TEST: c07s03b05x00p14n01i02541 - Type conversion can only occur on operand of universal real or integer."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c07s03b05x00p14n01i02541arch;
