entity emptyrec is
  port (
    clk_i           : in  bit
  );
end emptyrec;

architecture arch of emptyrec is
  type t_counter_config is record
  end record;
begin
end arch;
