context is
library use T.context is