package p is
  constant c : natural := 1;

  --  Comment for :state_t:
  type state_t is (s1, s2, s3);
end p;
