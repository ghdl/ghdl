library ieee;
context ieee.ieee_std_context;

entity fifo is
  generic ( gen : integer := 8 );
end fifo;

architecture arch of fifo is begin end;

