
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc170.vhd,v 1.2 2001-10-26 16:30:12 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c04s03b03x01p03n01i00170ent IS
END c04s03b03x01p03n01i00170ent;

ARCHITECTURE c04s03b03x01p03n01i00170arch OF c04s03b03x01p03n01i00170ent IS
  type x is range 1 to 10;
  signal Addr : bit;
  alias SIGN1 : x is x; -- fails_here
  alias SIGN2 : bit is Addr;
BEGIN
  TESTING: PROCESS
  BEGIN
    assert FALSE
      report "***FAILED TEST:c04s03b03x01p03n01i00170 - The name referred to in the alias declaration for SIGN1 is not a static name that refers to an object."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c04s03b03x01p03n01i00170arch;
