library IEEE;
use     IEEE.std_logic_1164.all;

entity ex1_entity is
  port (
    X : inout std_logic
  );
end entity;

architecture a of ex1_entity is
begin
end architecture;
