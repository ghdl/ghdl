entity name2 is
end name2;

architecture behav of name2 is
  signal samples: bit;
begin
  process
  begin
    bit'samples);
  end process;
end behav;
