entity entity_1 is
end entity entity_1;

architecture behav of entity_1 is
begin
	genIf: if True generate
		constant G0 : boolean := False;
	begin

	elsif False generate
		constant G1 : boolean := False;
	begin

	else generate
		constant G2 : boolean := False;
	begin

	end generate;
end architecture behav;
