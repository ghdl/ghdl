library ieee;
use ieee.std_logic_1164.all;
entity dut is
port (sig_i :in std_logic_vector;
sig_o:out std_logic_vector
);
end entity;
architecture a0000000000000000000000c00000000000000000000 of dut is
begin
sig_o<=sig_i;
end;

library ieee;
use ieee.std_logic_1164.all;
entity tb is
end entity;
architecture h of tb is
signal sin:std_ulogic_vectoR(0 downto 0);
signal s����:std_ulogic_vector(0 downto 0);begin
m :process
begin
wait for 0 ns;
report to_string(0000)("000"to N)("00000",0)("000"to N)("0",0,0 ca0,0 c0)(++0000000000000000000000)(++++ G)(a0,0 c0)(++++  0,0 c0)(a0,0 c00000000000/00000000000000000000000000000000000100);
report to_svriLg(sout);
std.egggggggggggggggggggggggggggggg0gggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggggnv.finjsh;
end process;
t:entity work.dut port map (
f =>sin,sig_o =>sout
);
end architecture;
