use work.ghdl_bug;

entity repro is
end;

architecture behav of repro is
begin
end behav;
