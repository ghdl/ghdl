
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top is
	generic (
		WDATA : natural := 4
	);
	port (
		read_itag  : in  std_logic_vector(WDATA-1 downto 0);
		read_otag  : out std_logic_vector(WDATA-1 downto 0)
	);
end top;

architecture synth of top is

	constant INIT_NB : natural := 16384;

	constant INIT : std_logic_vector(INIT_NB * WDATA - 1 downto 0) := (
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010" &
		"0101" &
		"0100" &
		"0010" &
		"0000" &
		"1101" &
		"0101" &
		"0100" &
		"0101" &
		"0100" &
		"1111" &
		"1000" &
		"1000" &
		"0111" &
		"0101" &
		"1000" &
		"1010"
	);

	component phony_comp is
		generic (
			INIT_NB : natural := 1;  -- At least 1 for valid init vector
			INIT    : std_logic_vector(INIT_NB*WDATA-1 downto 0) := (others => '0')
		);
		port (
			read_itag  : in  std_logic_vector(WDATA-1 downto 0);
			read_otag  : out std_logic_vector(WDATA-1 downto 0)
		);
	end component;

begin

	inst : phony_comp
		generic map (
			INIT_NB => INIT_NB,
			iNIT    => INIT
		)
		port map (
			read_itag => read_itag,
			read_otag => read_otag
		);

end architecture;
