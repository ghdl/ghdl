
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2966.vhd,v 1.2 2001-10-26 16:29:50 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c02s03b01x00p01n01i02966ent IS
END c02s03b01x00p01n01i02966ent;

ARCHITECTURE c02s03b01x00p01n01i02966arch OF c02s03b01x00p01n01i02966ent IS

BEGIN
  TESTING: PROCESS
    function "and" (a, b: in integer) return boolean is
    begin
      return false;
    end;
    variable i1, i2    :integer := 2;
    variable b1, b2    :boolean := true;
    variable q1      :boolean ;
    variable q2      :boolean ;
    variable q3      :boolean ;
  BEGIN
    q1 := i1 and i2;
    q2 := b1 and b2;
    q3 := "and" (i1, i2);
    wait for 5 ns;
    assert NOT( q1=false and q2=true and q3=false )
      report "***PASSED TEST: c02s03b01x00p01n01i02966"
      severity NOTE;
    assert ( q1=false and q2=true and q3=false )
      report "***FAILED TEST: c02s03b01x00p01n01i02966 - Function overload test failed."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c02s03b01x00p01n01i02966arch;
