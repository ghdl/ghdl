entity a is
 begin
   if r0  use
     type s array (n000000 range <>, block, c0000_000000);
                                     end if;
   end;
