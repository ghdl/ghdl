package function""begin r';