package gen0 is
generic(v:natural:=0);function get return natural;end;package body gen0 is
function get return natural is begin return 0;end;end gen0;package n is generic(package g is new n generic map(<>));function t return l;end;package body gen0 is use d;end gen0;package g is new n;package p is
end;architecture behav of b is
begin end behav;