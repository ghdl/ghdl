
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2515.vhd,v 1.2 2001-10-26 16:29:48 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c07s03b05x00p03n02i02515ent IS
END c07s03b05x00p03n02i02515ent;

ARCHITECTURE c07s03b05x00p03n02i02515arch OF c07s03b05x00p03n02i02515ent IS

BEGIN
  TESTING: PROCESS
    type century is range 1 to 10;
    
    function f(a:century) return century is
    begin 
      return century'(1); 
    end;
    
    type millenia is ('1', '2', '3', '4', '5');
    
    function f (a:millenia) return millenia is
    begin 
      return millenia'('2'); 
    end;
    
    variable hundreds : century  ;
  BEGIN
    hundreds := century (f(hundreds));
    assert NOT(hundreds = 1) 
      report "***PASSED TEST: c07s03b05x00p03n02i02515" 
      severity NOTE;
    assert (hundreds = 1) 
      report "***FAILED TEST: c07s03b05x00p03n02i02515 - Type of operand must be determinable independent of the context."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c07s03b05x00p03n02i02515arch;
