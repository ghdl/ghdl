package function is;s';