
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc764.vhd,v 1.2 2001-10-26 16:30:27 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

package c01s01b01x02p04n06i00764pkg is
  type ar_sig_range    is range 1 to 8;
  type ar_signal    is array (ar_sig_range) of BIT;
end c01s01b01x02p04n06i00764pkg;

use WORK.c01s01b01x02p04n06i00764pkg.all;
ENTITY c01s01b01x02p04n06i00764ent IS
  port (iface_array : ar_signal;
        iface_index : ar_sig_range);
END c01s01b01x02p04n06i00764ent;

ARCHITECTURE c01s01b01x02p04n06i00764arch OF c01s01b01x02p04n06i00764ent IS
  component COM_1 
    port ( F1 : in BIT);
  end component;
BEGIN
  CIS1: COM_1 
    port map ( iface_array (iface_index)); -- Failure_here
  --  Signal must be denoted by a static name

  TESTING: PROCESS
  BEGIN
    assert FALSE 
      report "***FAILED TEST: c01s01b01x02p04n06i00764 - Associated actual does not have a static name."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c01s01b01x02p04n06i00764arch;
