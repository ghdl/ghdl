library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

package pack_1 is
	constant const_1 : boolean := false;

end package;

package body pack_1 is
	constant const_1 : boolean := true;

end package body;
