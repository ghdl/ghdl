
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc228.vhd,v 1.2 2001-10-26 16:29:46 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s01b01x00p07n01i00228ent IS
END c03s01b01x00p07n01i00228ent;

ARCHITECTURE c03s01b01x00p07n01i00228arch OF c03s01b01x00p07n01i00228ent IS
  type MVL is ('0', '1', 'Z') ;
  type MVL1 is ('0', '1', 'Z', 'X') ;
  signal S1 : MVL ;
BEGIN
  TESTING: PROCESS
  BEGIN
    S1 <= '1' after 10 ns,
          '0' after 20 ns,
          'Z' after 50 ns; 
    wait for 60 ns;
    assert NOT( S1 = 'Z' )
      report "***PASSED TEST: c03s01b01x00p07n01i00228"
      severity NOTE;
    assert ( S1 = 'Z' )
      report "***FAILED TEST: c03s01b01x00p07n01i00228 - The type of an overloaded enumeration literal is determinable from the context."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s01b01x00p07n01i00228arch;
