library mwe;

entity mwe is
end entity;

architecture a of mwe is
begin
  process
  begin
    wait;
  end process;
end;
