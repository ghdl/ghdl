configuration cfg2 of e2 is
  -- comments in design units (python doc-string style) :cfg2:
  -- might be multi line :cfg2:
  for a2
  end for;
end configuration;
