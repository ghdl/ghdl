architecture a2 of e2 is
  -- comments in design units (python doc-string style) :a2:
    --:a2: might be multi line
begin

end architecture;
