entity ent1 is
end entity;

architecture rtl of ent1 is
 signal bwe : bit_vector (3 downto 0);
begin
end architecture;
