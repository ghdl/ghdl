library ieee;
use ieee.numeric_std.all;

package MyPkg is

  alias BCDType is unsigned(3 downto 0);

end package MyPkg;
