package pkg is
  type enum_t is (alpha, beta);
  alias alias_t is enum_t;
end package;

