entity tester is
end entity;

architecture a of tester is
    component check is
    end component;
begin
    checker: check;
end architecture;
