
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1014.vhd,v 1.2 2001-10-26 16:30:05 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c06s03b00x00p10n01i01014ent IS
END c06s03b00x00p10n01i01014ent;

ARCHITECTURE c06s03b00x00p10n01i01014arch OF c06s03b00x00p10n01i01014ent IS
  signal p : bit := '0';
  signal q : bit := '1';
BEGIN
  TESTING: PROCESS(c06s03b00x00p10n01i01014arch.p,c06s03b00x00p10n01i01014ent.q)
  BEGIN
    c06s03b00x00p10n01i01014ent.q <= c06s03b00x00p10n01i01014arch.p;
    assert FALSE 
      report "***FAILED TEST: c06s03b00x00p10n01i01014 - Declaration of suffix must occur within the construct denoted by the prefix."
      severity ERROR;
  END PROCESS TESTING;

END c06s03b00x00p10n01i01014arch;
