
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1436.vhd,v 1.2 2001-10-26 16:30:10 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c08s07b00x00p02n01i01436ent IS
END c08s07b00x00p02n01i01436ent;

ARCHITECTURE c08s07b00x00p02n01i01436arch OF c08s07b00x00p02n01i01436ent IS
begin

  TEST_PROCESS:  process
    variable I : INTEGER := 47;
  begin
    -- 'else' before 'elsif'.
    if  (I /= 47) then
      NULL;
    else
      NULL;
    elsif (I = 47) then
      NULL;
    end if;
    assert FALSE 
      report "***FAILED TEST: c08s07b00x00p02n01i01436 - reserved word 'elsif' is misplaced"
      severity ERROR;
    wait;
  end process TEST_PROCESS;

END c08s07b00x00p02n01i01436arch;
