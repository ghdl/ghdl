
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc3019.vhd,v 1.2 2001-10-26 16:30:24 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

package body c11s02b00x00p14n01i03019pkg is                   --- Failure_here
  type MVL2 is ('0','1','X','Z') ;
end c11s02b00x00p14n01i03019pkg;

ENTITY c11s02b00x00p14n01i03019ent IS
END c11s02b00x00p14n01i03019ent;

ARCHITECTURE c11s02b00x00p14n01i03019arch OF c11s02b00x00p14n01i03019ent IS

BEGIN
  TESTING: PROCESS
  BEGIN
    assert FALSE
      report "***FAILED TEST: c11s02b00x00p14n01i03019 - Secondary unit must reside in the same library as the primary unit."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c11s02b00x00p14n01i03019arch;
