library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ent is
end entity ent;

architecture arch of ent is
  signal test: natural;
begin
  LL: case test generate
    when =>
  end generate;
end architecture arch;
