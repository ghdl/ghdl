
architecture rtl of unit_b is
begin

    b <= not a;

end architecture;
