entity e is
end entity;

architecture a of e is
begin
end architecture;

