entity e is end entity;
architecture f of e is
signal foo: bit;
signal bar: bit;
begin
foo <= '1';
bar <= '0';
end f;
