entity test is
type type_test is range 0 to 2#1.1#2; -- here is the missing e between 2nd hash and 2
end;

