package p is
  --  Comment for the decl :c1:
  constant c1 : natural := 3;
end p;
