package phys is
type ANGLE is range INTEGER'range units
  sec;
  min = 60 sec;
  deg = 60 min;
end units;
end phys;
