
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc3056.vhd,v 1.2 2001-10-26 16:30:30 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

package c12s03b01x00p02n03i03056pkg is
  subtype BYTE is BIT_VECTOR(7 downto 0);
  function BIN_TO_INTG (IN_DATA : BYTE) return INTEGER;
end c12s03b01x00p02n03i03056pkg;

use WORK.c12s03b01x00p02n03i03056pkg.all;
ENTITY c12s03b01x00p02n03i03056ent IS
END c12s03b01x00p02n03i03056ent;

ARCHITECTURE c12s03b01x00p02n03i03056arch OF c12s03b01x00p02n03i03056ent IS

BEGIN
  TESTING: PROCESS
    variable S1 : BYTE := "00001111";
    variable X  : INTEGER;
  BEGIN
    X := BIN_TO_INTG(S1) ;
    assert FALSE
      report "***FAILED TEST: c12s03b01x00p02n03i03056 - Subprogram Body should be elaaborated before subprogram call."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c12s03b01x00p02n03i03056arch;
