-- comments before design units (javadoc / .net documentation style) :e1:
-- might be multiline :e1:
entity e1 is
end entity;
