architecture;l';