
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc313.vhd,v 1.2 2001-10-26 16:29:51 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s01b04x01p01n02i00313ent IS
END c03s01b04x01p01n02i00313ent;

ARCHITECTURE c03s01b04x01p01n02i00313arch OF c03s01b04x01p01n02i00313ent IS
  constant C1 : REAL := -1.0E38 ;
  constant C2 : REAL := +1.0E38 ;
BEGIN
  TESTING: PROCESS
    variable k1 : real;
    variable k2 : real;
  BEGIN
    k1 := C1;
    k2 := C2;
    assert NOT(k1=C1 and k2=C2)
      report "***PASSED TEST: c03s01b04x01p01n02i00313"
      severity NOTE;
    assert (k1=C1 and k2=C2)
      report "***FAILED TEST: c03s01b04x01p01n02i00313 - The range of REAL is host-independent, but it is guaranteed to include the range -1E38 to +1E38."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s01b04x01p01n02i00313arch;
