entity bug3 is
end;

architecture behavior of bug3 is
begin
    name(1 downto 0);
end behavior;
