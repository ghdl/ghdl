architecture if''h';