package pkg is
  constant cst : natural := 5;
end pkg;
