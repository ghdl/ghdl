
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc3017.vhd,v 1.2 2001-10-26 16:30:24 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

library lib01;
use lib01.c11s02b00x00p05n03i03017pkg.all;

ENTITY c11s02b00x00p05n03i03017ent IS
  assert my_bool
    report "Library clause preceeding entity is valid in entity scope."
    severity note;
END c11s02b00x00p05n03i03017ent;


use lib01.c11s02b00x00p05n03i03017pkg.all;         -- lib01 unknown Failed_here
ENTITY c11s02b00x00p05n03i03017ent IS
  assert my_bool
    report "Library clause is valid outside entity scope - test fails."
    severity note ;
END c11s02b00x00p05n03i03017ent;

ARCHITECTURE c11s02b00x00p05n03i03017arch OF c11s02b00x00p05n03i03017ent IS

BEGIN
  TESTING: PROCESS
  BEGIN
    assert FALSE
      report "***FAILED TEST: c11s02b00x00p05n03i03017 - Library clause only extends to the end of the declatative region associated with the design unit"
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c11s02b00x00p05n03i03017arch;
