library IEEE;
context IEEE.IEEE_std_context;

package my_fixed_pkg is new IEEE.fixed_generic_pkg;

--!

