architecture arch of ent is
  --  Comment
  signal b2 : bit;
begin
end arch;
