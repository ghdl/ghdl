package pkg2 is new work.gen2 generic map (work.pkg1);
