
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc283.vhd,v 1.2 2001-10-26 16:30:23 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s01b03x00p10n01i00283ent IS
END c03s01b03x00p10n01i00283ent;

ARCHITECTURE c03s01b03x00p10n01i00283arch OF c03s01b03x00p10n01i00283ent IS
  type J is               -- physical type decl
    range 0 to 1000
    units
      A;
      B = 10 A;
      C = 10.1 B;     -- Failure_here
      D = 10 C;
    end units;
BEGIN
  TESTING: PROCESS
  BEGIN
    assert FALSE 
      report "***FAILED TEST: c03s01b03x00p10n01i00283 - Abstract literal portion of a physical literal appearing in a secondary unit declaration must be integer literal."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s01b03x00p10n01i00283arch;
