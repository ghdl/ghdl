package pkga is
  subtype word is bit_vector (0 to 31);
end pkga;

