D%