entity repro2 is
end;

architecture behav of repro2 is
begin
   process
   begin
    "and";
   end process;
end;
