library ieee;
use ieee.std_logic_1164.all;

library ieee;
use ieee.numeric_std.all;

entity fsm_163 is
	port (
		clock : in  std_logic;
		reset : in  std_logic;
		out91 : out std_logic;
		out92 : out std_logic;
		out93 : out std_logic;
		in7 : in  std_logic;
		out94 : out std_logic;
		out95 : out std_logic;
		out98 : out std_logic;
		out100 : out std_logic;
		out101 : out std_logic;
		out102 : out std_logic;
		out104 : out std_logic;
		out105 : out std_logic;
		out106 : out std_logic;
		out107 : out std_logic;
		out108 : out std_logic;
		out109 : out std_logic;
		out111 : out std_logic;
		out114 : out std_logic;
		out116 : out std_logic;
		out118 : out std_logic;
		out119 : out std_logic;
		out120 : out std_logic;
		out128 : out std_logic;
		out130 : out std_logic;
		out131 : out std_logic;
		out132 : out std_logic;
		out137 : out std_logic;
		in8 : in  std_logic;
		out152 : out std_logic;
		out155 : out std_logic;
		out156 : out std_logic;
		out31 : out std_logic;
		in2 : in  std_logic;
		out28 : out std_logic;
		out29 : out std_logic;
		out30 : out std_logic;
		out26 : out std_logic;
		out27 : out std_logic;
		out24 : out std_logic;
		out25 : out std_logic;
		out77 : out std_logic;
		out79 : out std_logic;
		out80 : out std_logic;
		out82 : out std_logic;
		out34 : out std_logic;
		out35 : out std_logic;
		out36 : out std_logic;
		out32 : out std_logic;
		out33 : out std_logic;
		out40 : out std_logic;
		out41 : out std_logic;
		out88 : out std_logic;
		out89 : out std_logic;
		out21 : out std_logic;
		out22 : out std_logic;
		out23 : out std_logic;
		out73 : out std_logic;
		out76 : out std_logic;
		in6 : in  std_logic;
		out70 : out std_logic;
		out12 : out std_logic;
		out13 : out std_logic;
		out14 : out std_logic;
		out17 : out std_logic;
		out18 : out std_logic;
		out19 : out std_logic;
		out20 : out std_logic;
		out9 : out std_logic;
		out11 : out std_logic;
		out8 : out std_logic;
		out2 : out std_logic;
		out4 : out std_logic;
		out5 : out std_logic;
		in1 : in  std_logic;
		out6 : out std_logic;
		out7 : out std_logic;
		out0 : out std_logic;
		out1 : out std_logic;
		out37 : out std_logic;
		out38 : out std_logic;
		out39 : out std_logic;
		out1222 : out std_logic;
		out1223 : out std_logic;
		out1224 : out std_logic;
		out1225 : out std_logic;
		out1226 : out std_logic;
		out1228 : out std_logic;
		out1230 : out std_logic;
		in0 : in  std_logic;
		out67 : out std_logic;
		out68 : out std_logic;
		out65 : out std_logic;
		out66 : out std_logic;
		in5 : in  std_logic;
		out62 : out std_logic;
		out58 : out std_logic;
		out56 : out std_logic;
		in4 : in  std_logic;
		out57 : out std_logic;
		out54 : out std_logic;
		out55 : out std_logic;
		out51 : out std_logic;
		out52 : out std_logic;
		out53 : out std_logic;
		in3 : in  std_logic;
		out46 : out std_logic;
		out47 : out std_logic;
		out48 : out std_logic;
		out49 : out std_logic;
		out50 : out std_logic;
		out42 : out std_logic;
		out43 : out std_logic;
		out44 : out std_logic;
		out45 : out std_logic;
		in9 : in  std_logic;
		in10 : in  std_logic;
		out171 : out std_logic;
		in11 : in  std_logic;
		out191 : out std_logic;
		out207 : out std_logic;
		out208 : out std_logic;
		out209 : out std_logic;
		out212 : out std_logic;
		out213 : out std_logic;
		out216 : out std_logic;
		out220 : out std_logic;
		out221 : out std_logic;
		out223 : out std_logic;
		out224 : out std_logic;
		out226 : out std_logic;
		out227 : out std_logic;
		out228 : out std_logic;
		out229 : out std_logic;
		out230 : out std_logic;
		out233 : out std_logic;
		out235 : out std_logic;
		out236 : out std_logic;
		out237 : out std_logic;
		out238 : out std_logic;
		out239 : out std_logic;
		out241 : out std_logic;
		out250 : out std_logic;
		out258 : out std_logic;
		out259 : out std_logic;
		out261 : out std_logic;
		out270 : out std_logic;
		out276 : out std_logic;
		out277 : out std_logic;
		out283 : out std_logic;
		out285 : out std_logic;
		out287 : out std_logic;
		out290 : out std_logic;
		out291 : out std_logic;
		out293 : out std_logic;
		out301 : out std_logic;
		out303 : out std_logic;
		out304 : out std_logic;
		out315 : out std_logic;
		out319 : out std_logic;
		out321 : out std_logic;
		out330 : out std_logic;
		out335 : out std_logic;
		out338 : out std_logic;
		out341 : out std_logic;
		out342 : out std_logic;
		out344 : out std_logic;
		out347 : out std_logic;
		out351 : out std_logic;
		out354 : out std_logic;
		out355 : out std_logic;
		out356 : out std_logic;
		out357 : out std_logic;
		out358 : out std_logic;
		out360 : out std_logic;
		out361 : out std_logic;
		out362 : out std_logic;
		out365 : out std_logic;
		out367 : out std_logic;
		out368 : out std_logic;
		out370 : out std_logic;
		out375 : out std_logic;
		out376 : out std_logic;
		out378 : out std_logic;
		out381 : out std_logic;
		out382 : out std_logic;
		out386 : out std_logic;
		out387 : out std_logic;
		out388 : out std_logic;
		out390 : out std_logic;
		out392 : out std_logic;
		out393 : out std_logic;
		out394 : out std_logic;
		out397 : out std_logic;
		out403 : out std_logic;
		out404 : out std_logic;
		out408 : out std_logic;
		out409 : out std_logic;
		out410 : out std_logic;
		out412 : out std_logic;
		out416 : out std_logic;
		out417 : out std_logic;
		out418 : out std_logic;
		out419 : out std_logic;
		out420 : out std_logic;
		out421 : out std_logic;
		out424 : out std_logic;
		out425 : out std_logic;
		out430 : out std_logic;
		out431 : out std_logic;
		out434 : out std_logic;
		out436 : out std_logic;
		out438 : out std_logic;
		out439 : out std_logic;
		out440 : out std_logic;
		out441 : out std_logic;
		out442 : out std_logic;
		out443 : out std_logic;
		out444 : out std_logic;
		out445 : out std_logic;
		out446 : out std_logic;
		out447 : out std_logic;
		out448 : out std_logic;
		out450 : out std_logic;
		out451 : out std_logic;
		out454 : out std_logic;
		out457 : out std_logic;
		out460 : out std_logic;
		out463 : out std_logic;
		out465 : out std_logic;
		out466 : out std_logic;
		out472 : out std_logic;
		out473 : out std_logic;
		out475 : out std_logic;
		out476 : out std_logic;
		out479 : out std_logic;
		out480 : out std_logic;
		out481 : out std_logic;
		out482 : out std_logic;
		out484 : out std_logic;
		out485 : out std_logic;
		out489 : out std_logic;
		out491 : out std_logic;
		out494 : out std_logic;
		out497 : out std_logic;
		out500 : out std_logic;
		out503 : out std_logic;
		out504 : out std_logic;
		out505 : out std_logic;
		out508 : out std_logic;
		out509 : out std_logic;
		out513 : out std_logic;
		out514 : out std_logic;
		out516 : out std_logic;
		out521 : out std_logic;
		out523 : out std_logic;
		out524 : out std_logic;
		out525 : out std_logic;
		out530 : out std_logic;
		out532 : out std_logic;
		out533 : out std_logic;
		out535 : out std_logic;
		out536 : out std_logic;
		out539 : out std_logic;
		out541 : out std_logic;
		out543 : out std_logic;
		out545 : out std_logic;
		out547 : out std_logic;
		out549 : out std_logic;
		out550 : out std_logic;
		out552 : out std_logic;
		out558 : out std_logic;
		out559 : out std_logic;
		out563 : out std_logic;
		out566 : out std_logic;
		out572 : out std_logic;
		out573 : out std_logic;
		out576 : out std_logic;
		out577 : out std_logic;
		out581 : out std_logic;
		out582 : out std_logic;
		out590 : out std_logic;
		out591 : out std_logic;
		out592 : out std_logic;
		out593 : out std_logic;
		out595 : out std_logic;
		out611 : out std_logic;
		out619 : out std_logic;
		out638 : out std_logic;
		out643 : out std_logic;
		out644 : out std_logic;
		out645 : out std_logic;
		out646 : out std_logic;
		out648 : out std_logic;
		out650 : out std_logic;
		out652 : out std_logic;
		out657 : out std_logic;
		out659 : out std_logic;
		out662 : out std_logic;
		out677 : out std_logic;
		out678 : out std_logic;
		out679 : out std_logic;
		out680 : out std_logic;
		out682 : out std_logic;
		out686 : out std_logic;
		out692 : out std_logic;
		out1218 : out std_logic;
		out1219 : out std_logic;
		out1220 : out std_logic;
		out1221 : out std_logic;
		out695 : out std_logic;
		out697 : out std_logic;
		out706 : out std_logic;
		out719 : out std_logic;
		out729 : out std_logic;
		out744 : out std_logic;
		out746 : out std_logic;
		out748 : out std_logic;
		out833 : out std_logic;
		out834 : out std_logic;
		out836 : out std_logic;
		out837 : out std_logic;
		out839 : out std_logic;
		out840 : out std_logic;
		out841 : out std_logic;
		out844 : out std_logic;
		out845 : out std_logic;
		out846 : out std_logic;
		out848 : out std_logic;
		out850 : out std_logic;
		out852 : out std_logic;
		out854 : out std_logic;
		out856 : out std_logic;
		out858 : out std_logic;
		out860 : out std_logic;
		out863 : out std_logic;
		out865 : out std_logic;
		out866 : out std_logic;
		out873 : out std_logic;
		out877 : out std_logic;
		out888 : out std_logic;
		out891 : out std_logic;
		out893 : out std_logic;
		out895 : out std_logic;
		out898 : out std_logic;
		out900 : out std_logic;
		out902 : out std_logic;
		out903 : out std_logic;
		out904 : out std_logic;
		out905 : out std_logic;
		out906 : out std_logic;
		out907 : out std_logic;
		out908 : out std_logic;
		out909 : out std_logic;
		out910 : out std_logic;
		out912 : out std_logic;
		out913 : out std_logic;
		out914 : out std_logic;
		out915 : out std_logic;
		out917 : out std_logic;
		out920 : out std_logic;
		out921 : out std_logic;
		out924 : out std_logic;
		out934 : out std_logic;
		out935 : out std_logic;
		out937 : out std_logic;
		out938 : out std_logic;
		out940 : out std_logic;
		out943 : out std_logic;
		out945 : out std_logic;
		out957 : out std_logic;
		out958 : out std_logic;
		out962 : out std_logic;
		out968 : out std_logic;
		out972 : out std_logic;
		out973 : out std_logic;
		out974 : out std_logic;
		out975 : out std_logic;
		out976 : out std_logic;
		out980 : out std_logic;
		out986 : out std_logic;
		out988 : out std_logic;
		out989 : out std_logic;
		out990 : out std_logic;
		out1004 : out std_logic;
		out1008 : out std_logic;
		out999 : out std_logic;
		out1000 : out std_logic;
		out1002 : out std_logic;
		out1003 : out std_logic;
		out1050 : out std_logic;
		out1052 : out std_logic;
		out1053 : out std_logic;
		out1055 : out std_logic;
		out1056 : out std_logic;
		out1057 : out std_logic;
		out1059 : out std_logic;
		out1015 : out std_logic;
		out1025 : out std_logic;
		out1026 : out std_logic;
		out1038 : out std_logic;
		out1039 : out std_logic;
		out1042 : out std_logic;
		out1043 : out std_logic;
		out1046 : out std_logic;
		out1048 : out std_logic;
		out1061 : out std_logic;
		out1063 : out std_logic;
		out1064 : out std_logic;
		out1067 : out std_logic;
		out1068 : out std_logic;
		out1069 : out std_logic;
		out1071 : out std_logic;
		out1073 : out std_logic;
		out1076 : out std_logic;
		out1077 : out std_logic;
		out1078 : out std_logic;
		out1080 : out std_logic;
		out1081 : out std_logic;
		out1083 : out std_logic;
		out1085 : out std_logic;
		out1087 : out std_logic;
		out1089 : out std_logic;
		out1092 : out std_logic;
		out1096 : out std_logic;
		out1100 : out std_logic;
		out1103 : out std_logic;
		out1115 : out std_logic;
		out1122 : out std_logic;
		out1123 : out std_logic;
		out1127 : out std_logic;
		out1130 : out std_logic;
		out1133 : out std_logic;
		out1138 : out std_logic;
		out1139 : out std_logic;
		out1140 : out std_logic;
		out1141 : out std_logic;
		out1142 : out std_logic;
		out1143 : out std_logic;
		out1144 : out std_logic;
		out1145 : out std_logic;
		out1146 : out std_logic;
		out1147 : out std_logic;
		out1148 : out std_logic;
		out1149 : out std_logic;
		out1150 : out std_logic;
		out1151 : out std_logic;
		out1152 : out std_logic;
		out1153 : out std_logic;
		out1154 : out std_logic;
		out1155 : out std_logic;
		out1156 : out std_logic;
		out1157 : out std_logic;
		out1158 : out std_logic;
		out1159 : out std_logic;
		out1160 : out std_logic;
		out1161 : out std_logic;
		out1162 : out std_logic;
		out1163 : out std_logic;
		out1164 : out std_logic;
		out1165 : out std_logic;
		out1166 : out std_logic;
		out1167 : out std_logic;
		out1168 : out std_logic;
		out1169 : out std_logic;
		out1170 : out std_logic;
		out1171 : out std_logic;
		out1172 : out std_logic;
		out1173 : out std_logic;
		out1174 : out std_logic;
		out1175 : out std_logic;
		out1176 : out std_logic;
		out1177 : out std_logic;
		out1178 : out std_logic;
		out1179 : out std_logic;
		out1180 : out std_logic;
		out1181 : out std_logic;
		out1182 : out std_logic;
		out1183 : out std_logic;
		out1184 : out std_logic;
		out1185 : out std_logic;
		out1186 : out std_logic;
		out1187 : out std_logic;
		out1188 : out std_logic;
		out1189 : out std_logic;
		out1190 : out std_logic;
		out1191 : out std_logic;
		out1192 : out std_logic;
		out1193 : out std_logic;
		out1194 : out std_logic;
		out1195 : out std_logic;
		out1196 : out std_logic;
		out1197 : out std_logic;
		out1198 : out std_logic;
		out1199 : out std_logic;
		out1200 : out std_logic;
		out1201 : out std_logic;
		out1202 : out std_logic;
		out1203 : out std_logic;
		out1204 : out std_logic;
		out1205 : out std_logic;
		out1206 : out std_logic;
		out1207 : out std_logic;
		out1208 : out std_logic;
		out1209 : out std_logic;
		out1210 : out std_logic;
		out1211 : out std_logic;
		out1212 : out std_logic;
		out1213 : out std_logic;
		out1214 : out std_logic;
		out1215 : out std_logic;
		out1216 : out std_logic;
		out1217 : out std_logic
	);
end fsm_163;

architecture augh of fsm_163 is

	signal state_cur  : std_logic_vector(0 to 523) := (141 => '1', others => '0');
	signal state_next : std_logic_vector(0 to 523) := (141 => '1', others => '0');

	-- Buffers for outputs
	signal out386_buf : std_logic := '0';
	signal out386_bufn : std_logic;
	signal out404_buf : std_logic := '0';
	signal out404_bufn : std_logic;
	signal out457_buf : std_logic := '0';
	signal out457_bufn : std_logic;
	signal out841_buf : std_logic := '0';
	signal out841_bufn : std_logic;
	signal out276_buf : std_logic := '0';
	signal out276_bufn : std_logic;
	signal out67_buf : std_logic := '0';
	signal out67_bufn : std_logic;
	signal out239_buf : std_logic := '0';
	signal out239_bufn : std_logic;
	signal out259_buf : std_logic := '0';
	signal out259_bufn : std_logic;
	signal out416_buf : std_logic := '0';
	signal out416_bufn : std_logic;
	signal out646_buf : std_logic := '0';
	signal out646_bufn : std_logic;
	signal out485_buf : std_logic := '0';
	signal out485_bufn : std_logic;
	signal out935_buf : std_logic := '0';
	signal out935_bufn : std_logic;
	signal out463_buf : std_logic := '0';
	signal out463_bufn : std_logic;
	signal out120_buf : std_logic := '0';
	signal out120_bufn : std_logic;
	signal out293_buf : std_logic := '0';
	signal out293_bufn : std_logic;
	signal out216_buf : std_logic := '0';
	signal out216_bufn : std_logic;
	signal out319_buf : std_logic := '0';
	signal out319_bufn : std_logic;
	signal out230_buf : std_logic := '0';
	signal out230_bufn : std_logic;
	signal out1_buf : std_logic := '0';
	signal out1_bufn : std_logic;
	signal out93_buf : std_logic := '0';
	signal out93_bufn : std_logic;
	signal out89_buf : std_logic := '0';
	signal out89_bufn : std_logic;
	signal out539_buf : std_logic := '0';
	signal out539_bufn : std_logic;
	signal out62_buf : std_logic := '0';
	signal out62_bufn : std_logic;
	signal out856_buf : std_logic := '0';
	signal out856_bufn : std_logic;
	signal out451_buf : std_logic := '0';
	signal out451_bufn : std_logic;
	signal out287_buf : std_logic := '0';
	signal out287_bufn : std_logic;
	signal out315_buf : std_logic := '0';
	signal out315_bufn : std_logic;
	signal out536_buf : std_logic := '0';
	signal out536_bufn : std_logic;
	signal out209_buf : std_logic := '0';
	signal out209_bufn : std_logic;
	signal out221_buf : std_logic := '0';
	signal out221_bufn : std_logic;
	signal out283_buf : std_logic := '0';
	signal out283_bufn : std_logic;
	signal out368_buf : std_logic := '0';
	signal out368_bufn : std_logic;
	signal out516_buf : std_logic := '0';
	signal out516_bufn : std_logic;
	signal out393_buf : std_logic := '0';
	signal out393_bufn : std_logic;
	signal out1008_buf : std_logic := '0';
	signal out1008_bufn : std_logic;
	signal out392_buf : std_logic := '0';
	signal out392_bufn : std_logic;
	signal out261_buf : std_logic := '0';
	signal out261_bufn : std_logic;
	signal out559_buf : std_logic := '0';
	signal out559_bufn : std_logic;
	signal out543_buf : std_logic := '0';
	signal out543_bufn : std_logic;
	signal out895_buf : std_logic := '0';
	signal out895_bufn : std_logic;
	signal out82_buf : std_logic := '0';
	signal out82_bufn : std_logic;
	signal out220_buf : std_logic := '0';
	signal out220_bufn : std_logic;
	signal out95_buf : std_logic := '0';
	signal out95_bufn : std_logic;
	signal out943_buf : std_logic := '0';
	signal out943_bufn : std_logic;
	signal out465_buf : std_logic := '0';
	signal out465_bufn : std_logic;
	signal out238_buf : std_logic := '0';
	signal out238_bufn : std_logic;
	signal out1025_buf : std_logic := '0';
	signal out1025_bufn : std_logic;
	signal out132_buf : std_logic := '0';
	signal out132_bufn : std_logic;
	signal out79_buf : std_logic := '0';
	signal out79_bufn : std_logic;
	signal out500_buf : std_logic := '0';
	signal out500_bufn : std_logic;
	signal out65_buf : std_logic := '0';
	signal out65_bufn : std_logic;
	signal out111_buf : std_logic := '0';
	signal out111_bufn : std_logic;
	signal out420_buf : std_logic := '0';
	signal out420_bufn : std_logic;
	signal out1076_buf : std_logic := '0';
	signal out1076_bufn : std_logic;
	signal out101_buf : std_logic := '0';
	signal out101_bufn : std_logic;
	signal out106_buf : std_logic := '0';
	signal out106_bufn : std_logic;
	signal out68_buf : std_logic := '0';
	signal out68_bufn : std_logic;
	signal out1069_buf : std_logic := '0';
	signal out1069_bufn : std_logic;
	signal out77_buf : std_logic := '0';
	signal out77_bufn : std_logic;
	signal out102_buf : std_logic := '0';
	signal out102_bufn : std_logic;
	signal out394_buf : std_logic := '0';
	signal out394_bufn : std_logic;
	signal out342_buf : std_logic := '0';
	signal out342_bufn : std_logic;
	signal out104_buf : std_logic := '0';
	signal out104_bufn : std_logic;
	signal out361_buf : std_logic := '0';
	signal out361_bufn : std_logic;
	signal out116_buf : std_logic := '0';
	signal out116_bufn : std_logic;
	signal out595_buf : std_logic := '0';
	signal out595_bufn : std_logic;
	signal out1004_buf : std_logic := '0';
	signal out1004_bufn : std_logic;
	signal out227_buf : std_logic := '0';
	signal out227_bufn : std_logic;
	signal out109_buf : std_logic := '0';
	signal out109_bufn : std_logic;
	signal out619_buf : std_logic := '0';
	signal out619_bufn : std_logic;
	signal out410_buf : std_logic := '0';
	signal out410_bufn : std_logic;
	signal out989_buf : std_logic := '0';
	signal out989_bufn : std_logic;
	signal out431_buf : std_logic := '0';
	signal out431_bufn : std_logic;
	signal out938_buf : std_logic := '0';
	signal out938_bufn : std_logic;
	signal out525_buf : std_logic := '0';
	signal out525_bufn : std_logic;
	signal out73_buf : std_logic := '0';
	signal out73_bufn : std_logic;
	signal out837_buf : std_logic := '0';
	signal out837_bufn : std_logic;
	signal out860_buf : std_logic := '0';
	signal out860_bufn : std_logic;
	signal out228_buf : std_logic := '0';
	signal out228_bufn : std_logic;
	signal out421_buf : std_logic := '0';
	signal out421_bufn : std_logic;
	signal out409_buf : std_logic := '0';
	signal out409_bufn : std_logic;
	signal out473_buf : std_logic := '0';
	signal out473_bufn : std_logic;
	signal out509_buf : std_logic := '0';
	signal out509_bufn : std_logic;
	signal out94_buf : std_logic := '0';
	signal out94_bufn : std_logic;
	signal out1048_buf : std_logic := '0';
	signal out1048_bufn : std_logic;
	signal out98_buf : std_logic := '0';
	signal out98_bufn : std_logic;
	signal out945_buf : std_logic := '0';
	signal out945_bufn : std_logic;
	signal out156_buf : std_logic := '0';
	signal out156_bufn : std_logic;
	signal out152_buf : std_logic := '0';
	signal out152_bufn : std_logic;

	-- Retiming: counters
	signal rtmcounter0 :      unsigned(4 downto 0) := (others => '0');
	signal rtmcounter0_next : unsigned(4 downto 0);

	-- Retiming: Output of comparators
	signal rtmcmp92 : std_logic;
	signal rtmcmp128 : std_logic;
	signal rtmcmp276 : std_logic;
	signal rtmcmp290 : std_logic;

	-- Don't understand why these two function declarations are needed...
	function "/=" (L, R: std_logic) return std_logic is
	begin
		if L /= R then
			return '1';
		end if;
		return '0';
	end function;
	function "=" (L, R: std_logic) return std_logic is
	begin
		if L = R then
			return '1';
		end if;
		return '0';
	end function;

begin

	-- Sequential process
	-- Set the current state

	process (clock)
	begin
		if rising_edge(clock) then

			-- Next state
			state_cur <= state_next;
			-- Buffers for outputs
			out386_buf <= out386_bufn;
			out404_buf <= out404_bufn;
			out457_buf <= out457_bufn;
			out841_buf <= out841_bufn;
			out276_buf <= out276_bufn;
			out67_buf <= out67_bufn;
			out239_buf <= out239_bufn;
			out259_buf <= out259_bufn;
			out416_buf <= out416_bufn;
			out646_buf <= out646_bufn;
			out485_buf <= out485_bufn;
			out935_buf <= out935_bufn;
			out463_buf <= out463_bufn;
			out120_buf <= out120_bufn;
			out293_buf <= out293_bufn;
			out216_buf <= out216_bufn;
			out319_buf <= out319_bufn;
			out230_buf <= out230_bufn;
			out1_buf <= out1_bufn;
			out93_buf <= out93_bufn;
			out89_buf <= out89_bufn;
			out539_buf <= out539_bufn;
			out62_buf <= out62_bufn;
			out856_buf <= out856_bufn;
			out451_buf <= out451_bufn;
			out287_buf <= out287_bufn;
			out315_buf <= out315_bufn;
			out536_buf <= out536_bufn;
			out209_buf <= out209_bufn;
			out221_buf <= out221_bufn;
			out283_buf <= out283_bufn;
			out368_buf <= out368_bufn;
			out516_buf <= out516_bufn;
			out393_buf <= out393_bufn;
			out1008_buf <= out1008_bufn;
			out392_buf <= out392_bufn;
			out261_buf <= out261_bufn;
			out559_buf <= out559_bufn;
			out543_buf <= out543_bufn;
			out895_buf <= out895_bufn;
			out82_buf <= out82_bufn;
			out220_buf <= out220_bufn;
			out95_buf <= out95_bufn;
			out943_buf <= out943_bufn;
			out465_buf <= out465_bufn;
			out238_buf <= out238_bufn;
			out1025_buf <= out1025_bufn;
			out132_buf <= out132_bufn;
			out79_buf <= out79_bufn;
			out500_buf <= out500_bufn;
			out65_buf <= out65_bufn;
			out111_buf <= out111_bufn;
			out420_buf <= out420_bufn;
			out1076_buf <= out1076_bufn;
			out101_buf <= out101_bufn;
			out106_buf <= out106_bufn;
			out68_buf <= out68_bufn;
			out1069_buf <= out1069_bufn;
			out77_buf <= out77_bufn;
			out102_buf <= out102_bufn;
			out394_buf <= out394_bufn;
			out342_buf <= out342_bufn;
			out104_buf <= out104_bufn;
			out361_buf <= out361_bufn;
			out116_buf <= out116_bufn;
			out595_buf <= out595_bufn;
			out1004_buf <= out1004_bufn;
			out227_buf <= out227_bufn;
			out109_buf <= out109_bufn;
			out619_buf <= out619_bufn;
			out410_buf <= out410_bufn;
			out989_buf <= out989_bufn;
			out431_buf <= out431_bufn;
			out938_buf <= out938_bufn;
			out525_buf <= out525_bufn;
			out73_buf <= out73_bufn;
			out837_buf <= out837_bufn;
			out860_buf <= out860_bufn;
			out228_buf <= out228_bufn;
			out421_buf <= out421_bufn;
			out409_buf <= out409_bufn;
			out473_buf <= out473_bufn;
			out509_buf <= out509_bufn;
			out94_buf <= out94_bufn;
			out1048_buf <= out1048_bufn;
			out98_buf <= out98_bufn;
			out945_buf <= out945_bufn;
			out156_buf <= out156_bufn;
			out152_buf <= out152_bufn;
			-- Retiming: counters
			rtmcounter0 <= rtmcounter0_next;

		end if;
	end process;

	-- Retiming: the counters

	rtmcounter0_next <= rtmcounter0 + 1 when (reset /= '1') and (
		(state_cur(290) = '1' and rtmcmp290 = '0') or (state_cur(276) = '1' and rtmcmp276 = '0') or (state_cur(128) = '1' and rtmcmp128 = '0') or (state_cur(92) = '1' and rtmcmp92 = '0')
		) else (others => '0');

	-- Next state bits

	state_next(0) <= (reset /= '1') and ( ( state_cur(90) and not ( (NOT(in0)) = '1' ) ) );
	state_next(1) <= (reset /= '1') and ( ( state_cur(86) and not ( (NOT(in1)) = '1' ) ) );
	state_next(2) <= (reset /= '1') and ( ( state_cur(44) and not ( (NOT(in0)) = '1' ) ) );
	state_next(3) <= (reset /= '1') and ( ( state_cur(201) and not ( (NOT(in0)) = '1' ) ) );
	state_next(4) <= (reset /= '1') and ( ( state_cur(48) and not ( (NOT(in0)) = '1' ) ) );
	state_next(5) <= (reset /= '1') and ( ( state_cur(6) and not ( (NOT(in0)) = '1' ) ) );
	state_next(6) <= (reset /= '1') and ( state_cur(32) or ( state_cur(6) and (NOT(in0)) = '1' ) );
	state_next(7) <= (reset /= '1') and ( ( state_cur(207) and not ( (NOT(in0)) = '1' ) ) );
	state_next(8) <= (reset /= '1') and ( ( state_cur(17) and not ( (NOT(in0)) = '1' ) ) );
	state_next(9) <= (reset /= '1') and ( ( state_cur(13) and not ( (NOT(in0)) = '1' ) ) );
	state_next(10) <= (reset /= '1') and ( state_cur(221) or ( state_cur(10) and (NOT(in0)) = '1' ) );
	state_next(11) <= (reset /= '1') and ( state_cur(83) or ( state_cur(11) and (NOT(in1)) = '1' ) );
	state_next(12) <= (reset /= '1') and ( state_cur(23) or ( state_cur(12) and (NOT(in0)) = '1' ) );
	state_next(13) <= (reset /= '1') and ( state_cur(321) or ( state_cur(13) and (NOT(in0)) = '1' ) );
	state_next(14) <= (reset /= '1') and ( state_cur(251) or ( state_cur(14) and (NOT(in0)) = '1' ) );
	state_next(15) <= (reset /= '1') and ( ( state_cur(263) and not ( (NOT(in0)) = '1' ) ) );
	state_next(16) <= (reset /= '1') and ( ( state_cur(188) and not ( (NOT(in0)) = '1' ) ) );
	state_next(17) <= (reset /= '1') and ( ( state_cur(17) and (NOT(in0)) = '1' ) or state_cur(9) );
	state_next(18) <= (reset /= '1') and ( ( state_cur(239) and not ( (NOT(in0)) = '1' ) ) );
	state_next(19) <= (reset /= '1') and ( ( state_cur(14) and not ( (NOT(in0)) = '1' ) ) );
	state_next(20) <= (reset /= '1') and ( ( state_cur(27) and not ( (NOT(in0)) = '1' ) ) );
	state_next(21) <= (reset /= '1') and ( state_cur(22) or ( state_cur(21) and (NOT(in0)) = '1' ) );
	state_next(22) <= (reset /= '1') and ( ( state_cur(26) and not ( (NOT(in0)) = '1' ) ) );
	state_next(23) <= (reset /= '1') and ( ( state_cur(117) and not ( (NOT(in0)) = '1' ) ) );
	state_next(24) <= (reset /= '1') and ( state_cur(254) or ( state_cur(24) and (NOT(in0)) = '1' ) );
	state_next(25) <= (reset /= '1') and ( ( state_cur(320) and not ( (NOT(in0)) = '1' ) ) );
	state_next(26) <= (reset /= '1') and ( ( state_cur(26) and (NOT(in0)) = '1' ) or state_cur(25) );
	state_next(27) <= (reset /= '1') and ( state_cur(81) or ( state_cur(27) and (NOT(in0)) = '1' ) );
	state_next(28) <= (reset /= '1') and ( state_cur(261) or ( state_cur(28) and (NOT(in0)) = '1' ) );
	state_next(29) <= (reset /= '1') and ( state_cur(198) or ( state_cur(29) and (NOT(in1)) = '1' ) );
	state_next(30) <= (reset /= '1') and ( ( state_cur(324) and not ( (NOT(in0)) = '1' ) ) );
	state_next(31) <= (reset /= '1') and ( ( state_cur(33) and not ( (NOT(in0)) = '1' ) ) );
	state_next(32) <= (reset /= '1') and ( ( state_cur(259) and not ( (NOT(in0)) = '1' ) ) );
	state_next(33) <= (reset /= '1') and ( state_cur(267) or ( state_cur(33) and (NOT(in0)) = '1' ) );
	state_next(34) <= (reset /= '1') and ( ( state_cur(34) and (NOT(in0)) = '1' ) or state_cur(31) );
	state_next(35) <= (reset /= '1') and ( state_cur(36) or ( state_cur(35) and (NOT(in0)) = '1' ) );
	state_next(36) <= (reset /= '1') and ( ( state_cur(34) and not ( (NOT(in0)) = '1' ) ) );
	state_next(37) <= (reset /= '1') and ( state_cur(38) or ( state_cur(37) and (NOT(in0)) = '1' ) );
	state_next(38) <= (reset /= '1') and ( ( state_cur(35) and not ( (NOT(in0)) = '1' ) ) );
	state_next(39) <= (reset /= '1') and ( ( state_cur(323) and not ( (NOT(in0)) = '1' ) ) );
	state_next(40) <= (reset /= '1') and ( ( state_cur(285) and not ( (NOT(in0)) = '1' ) ) );
	state_next(41) <= (reset /= '1') and ( ( state_cur(41) and (NOT(in0)) = '1' ) or state_cur(8) );
	state_next(42) <= (reset /= '1') and ( state_cur(180) or ( state_cur(42) and (NOT(in1)) = '1' ) );
	state_next(43) <= (reset /= '1') and ( ( state_cur(41) and not ( (NOT(in0)) = '1' ) ) );
	state_next(44) <= (reset /= '1') and ( state_cur(66) or ( state_cur(44) and (NOT(in0)) = '1' ) );
	state_next(45) <= (reset /= '1') and ( ( state_cur(37) and not ( (NOT(in0)) = '1' ) ) );
	state_next(46) <= (reset /= '1') and ( ( state_cur(46) and (NOT(in0)) = '1' ) or state_cur(43) );
	state_next(47) <= (reset /= '1') and ( ( state_cur(46) and not ( (NOT(in0)) = '1' ) ) );
	state_next(48) <= (reset /= '1') and ( ( state_cur(48) and (NOT(in0)) = '1' ) or state_cur(40) );
	state_next(49) <= (reset /= '1') and ( ( state_cur(49) and (NOT(in0)) = '1' ) or state_cur(18) );
	state_next(50) <= (reset /= '1') and ( ( state_cur(50) and (NOT(in0)) = '1' ) or state_cur(47) );
	state_next(51) <= (reset /= '1') and ( state_cur(53) or ( state_cur(51) and (NOT(in0)) = '1' ) );
	state_next(52) <= (reset /= '1') and ( state_cur(56) or ( state_cur(52) and (NOT(in0)) = '1' ) );
	state_next(53) <= (reset /= '1') and ( ( state_cur(52) and not ( (NOT(in0)) = '1' ) ) );
	state_next(54) <= (reset /= '1') and ( ( state_cur(51) and not ( (NOT(in0)) = '1' ) ) );
	state_next(55) <= (reset /= '1') and ( ( state_cur(55) and (NOT(in0)) = '1' ) or state_cur(54) );
	state_next(56) <= (reset /= '1') and ( ( state_cur(21) and not ( (NOT(in0)) = '1' ) ) );
	state_next(57) <= (reset /= '1') and ( ( state_cur(104) and not ( (NOT(in0)) = '1' ) ) );
	state_next(58) <= (reset /= '1') and ( ( state_cur(12) and not ( (NOT(in0)) = '1' ) ) );
	state_next(59) <= (reset /= '1') and ( ( state_cur(61) and not ( (NOT(in0)) = '1' ) ) );
	state_next(60) <= (reset /= '1') and ( ( state_cur(246) and not ( (NOT(in0)) = '1' ) ) );
	state_next(61) <= (reset /= '1') and ( state_cur(260) or ( state_cur(61) and (NOT(in0)) = '1' ) );
	state_next(62) <= (reset /= '1') and ( ( state_cur(65) and not ( (NOT(in0)) = '1' ) ) );
	state_next(63) <= (reset /= '1') and ( ( state_cur(24) and not ( (NOT(in0)) = '1' ) ) );
	state_next(64) <= (reset /= '1') and ( state_cur(277) or ( state_cur(64) and (NOT(in0)) = '1' ) );
	state_next(65) <= (reset /= '1') and ( state_cur(329) or ( state_cur(65) and (NOT(in0)) = '1' ) );
	state_next(66) <= (reset /= '1') and ( ( state_cur(256) and not ( (NOT(in0)) = '1' ) ) );
	state_next(67) <= (reset /= '1') and ( ( state_cur(67) and (NOT(in0)) = '1' ) or state_cur(62) );
	state_next(68) <= (reset /= '1') and ( ( state_cur(68) and (NOT(in0)) = '1' ) or state_cur(60) );
	state_next(69) <= (reset /= '1') and ( ( state_cur(258) and not ( (NOT(in0)) = '1' ) ) );
	state_next(70) <= (reset /= '1') and ( ( state_cur(278) and not ( (NOT(in0)) = '1' ) ) );
	state_next(71) <= (reset /= '1') and ( ( state_cur(255) and not ( (NOT(in1)) = '1' ) ) );
	state_next(72) <= (reset /= '1') and ( state_cur(85) or ( state_cur(72) and (NOT(in1)) = '1' ) );
	state_next(73) <= (reset /= '1') and ( ( state_cur(106) and not ( (NOT(in1)) = '1' ) ) );
	state_next(74) <= (reset /= '1') and ( ( state_cur(297) and not ( (NOT(in0)) = '1' ) ) );
	state_next(75) <= (reset /= '1') and ( ( state_cur(75) and (NOT(in0)) = '1' ) or state_cur(57) );
	state_next(76) <= (reset /= '1') and ( ( state_cur(272) and not ( (NOT(in0)) = '1' ) ) );
	state_next(77) <= (reset /= '1') and ( state_cur(199) or ( state_cur(77) and (NOT(in0)) = '1' ) );
	state_next(78) <= (reset /= '1') and ( state_cur(115) or ( state_cur(78) and (NOT(in1)) = '1' ) );
	state_next(79) <= (reset /= '1') and ( ( state_cur(42) and not ( (NOT(in1)) = '1' ) ) );
	state_next(80) <= (reset /= '1') and ( ( state_cur(80) and (NOT(in0)) = '1' ) or state_cur(7) );
	state_next(81) <= (reset /= '1') and ( ( state_cur(80) and not ( (NOT(in0)) = '1' ) ) );
	state_next(82) <= (reset /= '1') and ( ( state_cur(217) and not ( (NOT(in0)) = '1' ) ) );
	state_next(83) <= (reset /= '1') and ( ( state_cur(72) and not ( (NOT(in1)) = '1' ) ) );
	state_next(84) <= (reset /= '1') and ( ( state_cur(84) and (NOT(in0)) = '1' ) or state_cur(82) );
	state_next(85) <= (reset /= '1') and ( ( state_cur(29) and not ( (NOT(in1)) = '1' ) ) );
	state_next(86) <= (reset /= '1') and ( state_cur(195) or ( state_cur(86) and (NOT(in1)) = '1' ) );
	state_next(87) <= (reset /= '1') and ( ( state_cur(87) and (NOT(in0)) = '1' ) or state_cur(20) );
	state_next(88) <= (reset /= '1') and ( ( state_cur(288) and not ( (NOT(in0)) = '1' ) ) );
	state_next(89) <= (reset /= '1') and ( ( state_cur(140) and not ( (NOT(in0)) = '1' ) ) );
	state_next(90) <= (reset /= '1') and ( ( state_cur(90) and (NOT(in0)) = '1' ) or state_cur(89) );
	state_next(91) <= (reset /= '1') and ( state_cur(337) );
	state_next(92) <= (reset /= '1') and ( (state_cur(92) = '1' and rtmcmp92 = '0') or state_cur(336) );
	state_next(93) <= (reset /= '1') and ( state_cur(339) );
	state_next(94) <= (reset /= '1') and ( ( state_cur(175) and not ( (in4) = '1' ) ) );
	state_next(95) <= (reset /= '1') and ( state_cur(334) );
	state_next(96) <= (reset /= '1') and ( state_cur(333) );
	state_next(97) <= (reset /= '1') and ( state_cur(244) or ( state_cur(97) and (NOT(in0)) = '1' ) );
	state_next(98) <= (reset /= '1') and ( state_cur(228) );
	state_next(99) <= (reset /= '1') and ( state_cur(273) or state_cur(105) );
	state_next(100) <= (reset /= '1') and ( state_cur(203) );
	state_next(101) <= (reset /= '1') and ( ( state_cur(101) and (NOT(in0)) = '1' ) or state_cur(5) );
	state_next(102) <= (reset /= '1') and ( state_cur(98) );
	state_next(103) <= (reset /= '1') and ( state_cur(200) );
	state_next(104) <= (reset /= '1') and ( state_cur(111) or ( state_cur(104) and (NOT(in0)) = '1' ) );
	state_next(105) <= (reset /= '1') and ( state_cur(301) );
	state_next(106) <= (reset /= '1') and ( state_cur(214) or ( state_cur(106) and (NOT(in1)) = '1' ) );
	state_next(107) <= (reset /= '1') and ( rtmcmp276 );
	state_next(108) <= (reset /= '1') and ( state_cur(224) );
	state_next(109) <= (reset /= '1') and ( ( state_cur(310) and (in9) = '1' ) );
	state_next(110) <= (reset /= '1') and ( state_cur(222) or ( state_cur(110) and (NOT(in1)) = '1' ) );
	state_next(111) <= (reset /= '1') and ( ( state_cur(112) and not ( (NOT(in0)) = '1' ) ) );
	state_next(112) <= (reset /= '1') and ( state_cur(293) or ( state_cur(112) and (NOT(in0)) = '1' ) );
	state_next(113) <= (reset /= '1') and ( ( state_cur(304) and not ( (NOT(in0)) = '1' ) ) );
	state_next(114) <= (reset /= '1') and ( state_cur(523) or state_cur(129) );
	state_next(115) <= (reset /= '1') and ( ( state_cur(110) and not ( (NOT(in1)) = '1' ) ) );
	state_next(116) <= (reset /= '1') and ( state_cur(327) or ( state_cur(116) and (NOT(in0)) = '1' ) );
	state_next(117) <= (reset /= '1') and ( ( state_cur(117) and (NOT(in0)) = '1' ) or state_cur(2) );
	state_next(118) <= (reset /= '1') and ( state_cur(181) or ( state_cur(118) and (NOT(in0)) = '1' ) );
	state_next(119) <= (reset /= '1') and ( state_cur(274) );
	state_next(120) <= (reset /= '1') and ( ( state_cur(120) and (NOT(in0)) = '1' ) or state_cur(15) );
	state_next(121) <= (reset /= '1') and ( state_cur(227) or ( state_cur(121) and (NOT(in0)) = '1' ) );
	state_next(122) <= (reset /= '1') and ( ( state_cur(122) and (NOT(in0)) = '1' ) or state_cur(4) );
	state_next(123) <= (reset /= '1') and ( state_cur(303) );
	state_next(124) <= (reset /= '1') and ( state_cur(133) or ( state_cur(124) and (NOT(in0)) = '1' ) );
	state_next(125) <= (reset /= '1') and ( ( state_cur(343) and not ( (NOT(in1)) = '1' ) ) );
	state_next(126) <= (reset /= '1') and ( ( state_cur(314) and not ( (NOT(in0)) = '1' ) ) );
	state_next(127) <= (reset /= '1') and ( ( state_cur(127) and (NOT(in0)) = '1' ) or state_cur(126) );
	state_next(128) <= (reset /= '1') and ( (state_cur(128) = '1' and rtmcmp128 = '0') or state_cur(296) );
	state_next(129) <= (reset /= '1') and ( ( state_cur(208) and (in5) = '1' ) );
	state_next(130) <= (reset /= '1') and ( state_cur(137) or ( state_cur(130) and (NOT(in0)) = '1' ) );
	state_next(131) <= (reset /= '1') and ( ( state_cur(127) and not ( (NOT(in0)) = '1' ) ) );
	state_next(132) <= (reset /= '1') and ( state_cur(191) );
	state_next(133) <= (reset /= '1') and ( ( state_cur(118) and not ( (NOT(in0)) = '1' ) ) );
	state_next(134) <= (reset /= '1') and ( state_cur(172) );
	state_next(135) <= (reset /= '1') and ( state_cur(284) or ( state_cur(135) and (NOT(in0)) = '1' ) );
	state_next(136) <= (reset /= '1') and ( state_cur(230) or ( state_cur(136) and (NOT(in0)) = '1' ) );
	state_next(137) <= (reset /= '1') and ( ( state_cur(116) and not ( (NOT(in0)) = '1' ) ) );
	state_next(138) <= (reset /= '1') and ( ( state_cur(175) and (in4) = '1' ) );
	state_next(139) <= (reset /= '1') and ( ( state_cur(101) and not ( (NOT(in0)) = '1' ) ) );
	state_next(140) <= (reset /= '1') and ( ( state_cur(140) and (NOT(in0)) = '1' ) or state_cur(139) );
	state_next(141) <= (reset = '1') or ( ( state_cur(141) and (NOT(in2)) = '1' ) );
	state_next(142) <= (reset /= '1') and ( state_cur(270) );
	state_next(143) <= (reset /= '1') and ( state_cur(204) );
	state_next(144) <= (reset /= '1') and ( state_cur(173) );
	state_next(145) <= (reset /= '1') and ( state_cur(322) );
	state_next(146) <= (reset /= '1') and ( state_cur(331) );
	state_next(147) <= (reset /= '1') and ( state_cur(197) );
	state_next(148) <= (reset /= '1') and ( state_cur(306) );
	state_next(149) <= (reset /= '1') and ( state_cur(187) );
	state_next(150) <= (reset /= '1') and ( state_cur(294) );
	state_next(151) <= (reset /= '1') and ( state_cur(289) );
	state_next(152) <= (reset /= '1') and ( ( state_cur(153) and not ( (NOT(in0)) = '1' ) ) );
	state_next(153) <= (reset /= '1') and ( state_cur(154) or ( state_cur(153) and (NOT(in0)) = '1' ) );
	state_next(154) <= (reset /= '1') and ( ( state_cur(155) and not ( (NOT(in0)) = '1' ) ) );
	state_next(155) <= (reset /= '1') and ( state_cur(156) or ( state_cur(155) and (NOT(in0)) = '1' ) );
	state_next(156) <= (reset /= '1') and ( ( state_cur(157) and not ( (NOT(in0)) = '1' ) ) );
	state_next(157) <= (reset /= '1') and ( state_cur(158) or ( state_cur(157) and (NOT(in0)) = '1' ) );
	state_next(158) <= (reset /= '1') and ( ( state_cur(159) and not ( (NOT(in0)) = '1' ) ) );
	state_next(159) <= (reset /= '1') and ( state_cur(160) or ( state_cur(159) and (NOT(in0)) = '1' ) );
	state_next(160) <= (reset /= '1') and ( ( state_cur(161) and not ( (NOT(in0)) = '1' ) ) );
	state_next(161) <= (reset /= '1') and ( state_cur(162) or ( state_cur(161) and (NOT(in0)) = '1' ) );
	state_next(162) <= (reset /= '1') and ( ( state_cur(163) and not ( (NOT(in0)) = '1' ) ) );
	state_next(163) <= (reset /= '1') and ( state_cur(164) or ( state_cur(163) and (NOT(in0)) = '1' ) );
	state_next(164) <= (reset /= '1') and ( ( state_cur(165) and not ( (NOT(in0)) = '1' ) ) );
	state_next(165) <= (reset /= '1') and ( state_cur(166) or ( state_cur(165) and (NOT(in0)) = '1' ) );
	state_next(166) <= (reset /= '1') and ( ( state_cur(167) and not ( (NOT(in0)) = '1' ) ) );
	state_next(167) <= (reset /= '1') and ( state_cur(168) or ( state_cur(167) and (NOT(in0)) = '1' ) );
	state_next(168) <= (reset /= '1') and ( ( state_cur(55) and not ( (NOT(in0)) = '1' ) ) );
	state_next(169) <= (reset /= '1') and ( state_cur(332) );
	state_next(170) <= (reset /= '1') and ( state_cur(169) );
	state_next(171) <= (reset /= '1') and ( ( state_cur(171) and (NOT(in0)) = '1' ) or state_cur(16) );
	state_next(172) <= (reset /= '1') and ( state_cur(174) );
	state_next(173) <= (reset /= '1') and ( ( state_cur(325) and (in10) = '1' ) or ( state_cur(310) and not ( (in9) = '1' ) ) );
	state_next(174) <= (reset /= '1') and ( state_cur(319) );
	state_next(175) <= (reset /= '1') and ( state_cur(170) );
	state_next(176) <= (reset /= '1') and ( ( state_cur(176) and (NOT(in0)) = '1' ) or state_cur(70) );
	state_next(177) <= (reset /= '1') and ( ( state_cur(279) and not ( (NOT(in0)) = '1' ) ) );
	state_next(178) <= (reset /= '1') and ( ( state_cur(150) and (in3) = '1' ) );
	state_next(179) <= (reset /= '1') and ( state_cur(282) );
	state_next(180) <= (reset /= '1') and ( ( state_cur(520) and not ( (NOT(in1)) = '1' ) ) );
	state_next(181) <= (reset /= '1') and ( ( state_cur(226) and not ( (NOT(in0)) = '1' ) ) );
	state_next(182) <= (reset /= '1') and ( state_cur(223) );
	state_next(183) <= (reset /= '1') and ( state_cur(280) );
	state_next(184) <= (reset /= '1') and ( state_cur(183) );
	state_next(185) <= (reset /= '1') and ( ( state_cur(135) and not ( (NOT(in0)) = '1' ) ) );
	state_next(186) <= (reset /= '1') and ( rtmcmp290 );
	state_next(187) <= (reset /= '1') and ( state_cur(184) );
	state_next(188) <= (reset /= '1') and ( state_cur(206) or ( state_cur(188) and (NOT(in0)) = '1' ) );
	state_next(189) <= (reset /= '1') and ( state_cur(179) );
	state_next(190) <= (reset /= '1') and ( state_cur(186) );
	state_next(191) <= (reset /= '1') and ( state_cur(190) );
	state_next(192) <= (reset /= '1') and ( ( state_cur(192) and (NOT(in0)) = '1' ) or state_cur(76) );
	state_next(193) <= (reset /= '1') and ( state_cur(233) );
	state_next(194) <= (reset /= '1') and ( state_cur(252) or ( state_cur(194) and (NOT(in0)) = '1' ) );
	state_next(195) <= (reset /= '1') and ( ( state_cur(521) and not ( (NOT(in1)) = '1' ) ) );
	state_next(196) <= (reset /= '1') and ( state_cur(231) );
	state_next(197) <= (reset /= '1') and ( state_cur(218) );
	state_next(198) <= (reset /= '1') and ( ( state_cur(78) and not ( (NOT(in1)) = '1' ) ) );
	state_next(199) <= (reset /= '1') and ( ( state_cur(120) and not ( (NOT(in0)) = '1' ) ) );
	state_next(200) <= (reset /= '1') and ( state_cur(95) );
	state_next(201) <= (reset /= '1') and ( state_cur(307) or ( state_cur(201) and (NOT(in0)) = '1' ) );
	state_next(202) <= (reset /= '1') and ( state_cur(266) or ( state_cur(202) and (NOT(in0)) = '1' ) );
	state_next(203) <= (reset /= '1') and ( state_cur(91) );
	state_next(204) <= (reset /= '1') and ( state_cur(123) );
	state_next(205) <= (reset /= '1') and ( ( state_cur(211) and not ( (NOT(in0)) = '1' ) ) );
	state_next(206) <= (reset /= '1') and ( ( state_cur(136) and not ( (NOT(in0)) = '1' ) ) );
	state_next(207) <= (reset /= '1') and ( ( state_cur(207) and (NOT(in0)) = '1' ) or state_cur(205) );
	state_next(208) <= (reset /= '1') and ( state_cur(300) );
	state_next(209) <= (reset /= '1') and ( state_cur(312) );
	state_next(210) <= (reset /= '1') and ( state_cur(292) );
	state_next(211) <= (reset /= '1') and ( ( state_cur(211) and (NOT(in0)) = '1' ) or state_cur(185) );
	state_next(212) <= (reset /= '1') and ( state_cur(326) );
	state_next(213) <= (reset /= '1') and ( state_cur(340) );
	state_next(214) <= (reset /= '1') and ( ( state_cur(11) and not ( (NOT(in1)) = '1' ) ) );
	state_next(215) <= (reset /= '1') and ( state_cur(229) or ( state_cur(215) and (NOT(in0)) = '1' ) );
	state_next(216) <= (reset /= '1') and ( state_cur(248) or ( state_cur(216) and (NOT(in0)) = '1' ) );
	state_next(217) <= (reset /= '1') and ( state_cur(271) or ( state_cur(217) and (NOT(in0)) = '1' ) );
	state_next(218) <= (reset /= '1') and ( state_cur(146) or state_cur(138) );
	state_next(219) <= (reset /= '1') and ( state_cur(151) );
	state_next(220) <= (reset /= '1') and ( state_cur(298) );
	state_next(221) <= (reset /= '1') and ( ( state_cur(318) and not ( (NOT(in0)) = '1' ) ) );
	state_next(222) <= (reset /= '1') and ( state_cur(152) or ( state_cur(141) and not ( (NOT(in2)) = '1' ) ) );
	state_next(223) <= (reset /= '1') and ( state_cur(232) );
	state_next(224) <= (reset /= '1') and ( state_cur(342) );
	state_next(225) <= (reset /= '1') and ( ( state_cur(202) and not ( (NOT(in0)) = '1' ) ) );
	state_next(226) <= (reset /= '1') and ( state_cur(311) or ( state_cur(226) and (NOT(in0)) = '1' ) );
	state_next(227) <= (reset /= '1') and ( ( state_cur(250) and not ( (NOT(in0)) = '1' ) ) );
	state_next(228) <= (reset /= '1') and ( state_cur(189) );
	state_next(229) <= (reset /= '1') and ( ( state_cur(216) and not ( (NOT(in0)) = '1' ) ) );
	state_next(230) <= (reset /= '1') and ( ( state_cur(176) and not ( (NOT(in0)) = '1' ) ) );
	state_next(231) <= (reset /= '1') and ( state_cur(234) );
	state_next(232) <= (reset /= '1') and ( state_cur(145) );
	state_next(233) <= (reset /= '1') and ( state_cur(236) );
	state_next(234) <= (reset /= '1') and ( state_cur(235) );
	state_next(235) <= (reset /= '1') and ( state_cur(102) );
	state_next(236) <= (reset /= '1') and ( state_cur(237) );
	state_next(237) <= (reset /= '1') and ( state_cur(99) );
	state_next(238) <= (reset /= '1') and ( ( state_cur(287) and not ( (NOT(in0)) = '1' ) ) );
	state_next(239) <= (reset /= '1') and ( ( state_cur(239) and (NOT(in0)) = '1' ) or state_cur(58) );
	state_next(240) <= (reset /= '1') and ( state_cur(241) or state_cur(148) );
	state_next(241) <= (reset /= '1') and ( ( state_cur(245) and not ( (in8) = '1' ) ) );
	state_next(242) <= (reset /= '1') and ( ( state_cur(97) and not ( (NOT(in0)) = '1' ) ) );
	state_next(243) <= (reset /= '1') and ( state_cur(275) or ( state_cur(243) and (NOT(in0)) = '1' ) );
	state_next(244) <= (reset /= '1') and ( ( state_cur(245) and (in8) = '1' ) );
	state_next(245) <= (reset /= '1') and ( state_cur(247) or state_cur(242) );
	state_next(246) <= (reset /= '1') and ( state_cur(253) or ( state_cur(246) and (NOT(in0)) = '1' ) );
	state_next(247) <= (reset /= '1') and ( ( state_cur(328) and not ( (in11) = '1' ) ) );
	state_next(248) <= (reset /= '1') and ( ( state_cur(302) and not ( (NOT(in0)) = '1' ) ) );
	state_next(249) <= (reset /= '1') and ( ( state_cur(77) and not ( (NOT(in0)) = '1' ) ) );
	state_next(250) <= (reset /= '1') and ( ( state_cur(250) and (NOT(in0)) = '1' ) or state_cur(88) );
	state_next(251) <= (reset /= '1') and ( ( state_cur(130) and not ( (NOT(in0)) = '1' ) ) );
	state_next(252) <= (reset /= '1') and ( ( state_cur(171) and not ( (NOT(in0)) = '1' ) ) );
	state_next(253) <= (reset /= '1') and ( ( state_cur(49) and not ( (NOT(in0)) = '1' ) ) );
	state_next(254) <= (reset /= '1') and ( ( state_cur(68) and not ( (NOT(in0)) = '1' ) ) );
	state_next(255) <= (reset /= '1') and ( ( state_cur(255) and (NOT(in1)) = '1' ) or state_cur(79) );
	state_next(256) <= (reset /= '1') and ( ( state_cur(256) and (NOT(in0)) = '1' ) or state_cur(69) );
	state_next(257) <= (reset /= '1') and ( ( state_cur(64) and not ( (NOT(in0)) = '1' ) ) );
	state_next(258) <= (reset /= '1') and ( ( state_cur(258) and (NOT(in0)) = '1' ) or state_cur(249) );
	state_next(259) <= (reset /= '1') and ( state_cur(283) or ( state_cur(259) and (NOT(in0)) = '1' ) );
	state_next(260) <= (reset /= '1') and ( ( state_cur(50) and not ( (NOT(in0)) = '1' ) ) );
	state_next(261) <= (reset /= '1') and ( ( state_cur(269) and not ( (NOT(in0)) = '1' ) ) );
	state_next(262) <= (reset /= '1') and ( ( state_cur(240) and not ( (in7) = '1' ) ) );
	state_next(263) <= (reset /= '1') and ( ( state_cur(263) and (NOT(in0)) = '1' ) or state_cur(19) );
	state_next(264) <= (reset /= '1') and ( state_cur(315) or ( state_cur(264) and (NOT(in0)) = '1' ) );
	state_next(265) <= (reset /= '1') and ( ( state_cur(124) and not ( (NOT(in0)) = '1' ) ) );
	state_next(266) <= (reset /= '1') and ( ( state_cur(87) and not ( (NOT(in0)) = '1' ) ) );
	state_next(267) <= (reset /= '1') and ( ( state_cur(243) and not ( (NOT(in0)) = '1' ) ) );
	state_next(268) <= (reset /= '1') and ( state_cur(103) );
	state_next(269) <= (reset /= '1') and ( ( state_cur(269) and (NOT(in0)) = '1' ) or state_cur(257) );
	state_next(270) <= (reset /= '1') and ( state_cur(144) );
	state_next(271) <= (reset /= '1') and ( ( state_cur(28) and not ( (NOT(in0)) = '1' ) ) );
	state_next(272) <= (reset /= '1') and ( ( state_cur(272) and (NOT(in0)) = '1' ) or state_cur(225) );
	state_next(273) <= (reset /= '1') and ( ( state_cur(220) and (in6) = '1' ) );
	state_next(274) <= (reset /= '1') and ( state_cur(134) );
	state_next(275) <= (reset /= '1') and ( ( state_cur(75) and not ( (NOT(in0)) = '1' ) ) );
	state_next(276) <= (reset /= '1') and ( (state_cur(276) = '1' and rtmcmp276 = '0') or state_cur(114) );
	state_next(277) <= (reset /= '1') and ( ( state_cur(67) and not ( (NOT(in0)) = '1' ) ) );
	state_next(278) <= (reset /= '1') and ( ( state_cur(278) and (NOT(in0)) = '1' ) or state_cur(265) );
	state_next(279) <= (reset /= '1') and ( ( state_cur(279) and (NOT(in0)) = '1' ) or state_cur(3) );
	state_next(280) <= (reset /= '1') and ( state_cur(281) );
	state_next(281) <= (reset /= '1') and ( ( state_cur(208) and not ( (in5) = '1' ) ) );
	state_next(282) <= (reset /= '1') and ( state_cur(100) );
	state_next(283) <= (reset /= '1') and ( ( state_cur(10) and not ( (NOT(in0)) = '1' ) ) );
	state_next(284) <= (reset /= '1') and ( ( state_cur(264) and not ( (NOT(in0)) = '1' ) ) );
	state_next(285) <= (reset /= '1') and ( state_cur(286) or ( state_cur(285) and (NOT(in0)) = '1' ) );
	state_next(286) <= (reset /= '1') and ( ( state_cur(313) and not ( (NOT(in0)) = '1' ) ) );
	state_next(287) <= (reset /= '1') and ( ( state_cur(287) and (NOT(in0)) = '1' ) or state_cur(177) );
	state_next(288) <= (reset /= '1') and ( ( state_cur(288) and (NOT(in0)) = '1' ) or state_cur(45) );
	state_next(289) <= (reset /= '1') and ( state_cur(210) );
	state_next(290) <= (reset /= '1') and ( (state_cur(290) = '1' and rtmcmp290 = '0') or state_cur(291) );
	state_next(291) <= (reset /= '1') and ( ( state_cur(240) and (in7) = '1' ) );
	state_next(292) <= (reset /= '1') and ( state_cur(147) );
	state_next(293) <= (reset /= '1') and ( ( state_cur(295) and not ( (NOT(in0)) = '1' ) ) );
	state_next(294) <= (reset /= '1') and ( state_cur(132) );
	state_next(295) <= (reset /= '1') and ( ( state_cur(295) and (NOT(in0)) = '1' ) or state_cur(113) );
	state_next(296) <= (reset /= '1') and ( state_cur(268) or state_cur(178) );
	state_next(297) <= (reset /= '1') and ( ( state_cur(297) and (NOT(in0)) = '1' ) or state_cur(0) );
	state_next(298) <= (reset /= '1') and ( state_cur(143) );
	state_next(299) <= (reset /= '1') and ( ( state_cur(194) and not ( (NOT(in0)) = '1' ) ) );
	state_next(300) <= (reset /= '1') and ( state_cur(142) );
	state_next(301) <= (reset /= '1') and ( state_cur(108) );
	state_next(302) <= (reset /= '1') and ( ( state_cur(302) and (NOT(in0)) = '1' ) or state_cur(299) );
	state_next(303) <= (reset /= '1') and ( rtmcmp128 );
	state_next(304) <= (reset /= '1') and ( ( state_cur(304) and (NOT(in0)) = '1' ) or state_cur(39) );
	state_next(305) <= (reset /= '1') and ( ( state_cur(305) and (NOT(in0)) = '1' ) or state_cur(30) );
	state_next(306) <= (reset /= '1') and ( state_cur(209) );
	state_next(307) <= (reset /= '1') and ( ( state_cur(192) and not ( (NOT(in0)) = '1' ) ) );
	state_next(308) <= (reset /= '1') and ( ( state_cur(325) and not ( (in10) = '1' ) ) );
	state_next(309) <= (reset /= '1') and ( ( state_cur(122) and not ( (NOT(in0)) = '1' ) ) );
	state_next(310) <= (reset /= '1') and ( state_cur(308) or state_cur(196) );
	state_next(311) <= (reset /= '1') and ( ( state_cur(84) and not ( (NOT(in0)) = '1' ) ) );
	state_next(312) <= (reset /= '1') and ( state_cur(119) );
	state_next(313) <= (reset /= '1') and ( state_cur(330) or ( state_cur(313) and (NOT(in0)) = '1' ) );
	state_next(314) <= (reset /= '1') and ( ( state_cur(314) and (NOT(in0)) = '1' ) or state_cur(59) );
	state_next(315) <= (reset /= '1') and ( ( state_cur(121) and not ( (NOT(in0)) = '1' ) ) );
	state_next(316) <= (reset /= '1') and ( ( state_cur(316) and (NOT(in0)) = '1' ) or state_cur(63) );
	state_next(317) <= (reset /= '1') and ( ( state_cur(317) and (NOT(in0)) = '1' ) or state_cur(74) );
	state_next(318) <= (reset /= '1') and ( ( state_cur(318) and (NOT(in0)) = '1' ) or state_cur(262) );
	state_next(319) <= (reset /= '1') and ( state_cur(338) );
	state_next(320) <= (reset /= '1') and ( ( state_cur(320) and (NOT(in0)) = '1' ) or state_cur(131) );
	state_next(321) <= (reset /= '1') and ( ( state_cur(316) and not ( (NOT(in0)) = '1' ) ) );
	state_next(322) <= (reset /= '1') and ( state_cur(212) );
	state_next(323) <= (reset /= '1') and ( ( state_cur(323) and (NOT(in0)) = '1' ) or state_cur(309) );
	state_next(324) <= (reset /= '1') and ( ( state_cur(324) and (NOT(in0)) = '1' ) or state_cur(238) );
	state_next(325) <= (reset /= '1') and ( state_cur(109) );
	state_next(326) <= (reset /= '1') and ( state_cur(107) );
	state_next(327) <= (reset /= '1') and ( ( state_cur(215) and not ( (NOT(in0)) = '1' ) ) );
	state_next(328) <= (reset /= '1') and ( state_cur(219) or state_cur(125) );
	state_next(329) <= (reset /= '1') and ( ( state_cur(305) and not ( (NOT(in0)) = '1' ) ) );
	state_next(330) <= (reset /= '1') and ( ( state_cur(317) and not ( (NOT(in0)) = '1' ) ) );
	state_next(331) <= (reset /= '1') and ( state_cur(213) );
	state_next(332) <= (reset /= '1') and ( state_cur(335) );
	state_next(333) <= (reset /= '1') and ( ( state_cur(150) and not ( (in3) = '1' ) ) );
	state_next(334) <= (reset /= '1') and ( state_cur(96) );
	state_next(335) <= (reset /= '1') and ( state_cur(182) );
	state_next(336) <= (reset /= '1') and ( ( state_cur(328) and (in11) = '1' ) );
	state_next(337) <= (reset /= '1') and ( rtmcmp92 );
	state_next(338) <= (reset /= '1') and ( state_cur(193) );
	state_next(339) <= (reset /= '1') and ( state_cur(94) );
	state_next(340) <= (reset /= '1') and ( state_cur(93) );
	state_next(341) <= (reset /= '1') and ( state_cur(522) );
	state_next(342) <= (reset /= '1') and ( state_cur(341) );
	state_next(343) <= (reset /= '1') and ( state_cur(344) or ( state_cur(343) and (NOT(in1)) = '1' ) );
	state_next(344) <= (reset /= '1') and ( ( state_cur(345) and not ( (NOT(in1)) = '1' ) ) );
	state_next(345) <= (reset /= '1') and ( state_cur(346) or ( state_cur(345) and (NOT(in1)) = '1' ) );
	state_next(346) <= (reset /= '1') and ( ( state_cur(347) and not ( (NOT(in1)) = '1' ) ) );
	state_next(347) <= (reset /= '1') and ( state_cur(348) or ( state_cur(347) and (NOT(in1)) = '1' ) );
	state_next(348) <= (reset /= '1') and ( ( state_cur(349) and not ( (NOT(in1)) = '1' ) ) );
	state_next(349) <= (reset /= '1') and ( state_cur(350) or ( state_cur(349) and (NOT(in1)) = '1' ) );
	state_next(350) <= (reset /= '1') and ( ( state_cur(351) and not ( (NOT(in1)) = '1' ) ) );
	state_next(351) <= (reset /= '1') and ( state_cur(352) or ( state_cur(351) and (NOT(in1)) = '1' ) );
	state_next(352) <= (reset /= '1') and ( ( state_cur(353) and not ( (NOT(in1)) = '1' ) ) );
	state_next(353) <= (reset /= '1') and ( state_cur(354) or ( state_cur(353) and (NOT(in1)) = '1' ) );
	state_next(354) <= (reset /= '1') and ( ( state_cur(355) and not ( (NOT(in1)) = '1' ) ) );
	state_next(355) <= (reset /= '1') and ( state_cur(356) or ( state_cur(355) and (NOT(in1)) = '1' ) );
	state_next(356) <= (reset /= '1') and ( ( state_cur(357) and not ( (NOT(in1)) = '1' ) ) );
	state_next(357) <= (reset /= '1') and ( state_cur(358) or ( state_cur(357) and (NOT(in1)) = '1' ) );
	state_next(358) <= (reset /= '1') and ( ( state_cur(359) and not ( (NOT(in1)) = '1' ) ) );
	state_next(359) <= (reset /= '1') and ( state_cur(360) or ( state_cur(359) and (NOT(in1)) = '1' ) );
	state_next(360) <= (reset /= '1') and ( ( state_cur(361) and not ( (NOT(in1)) = '1' ) ) );
	state_next(361) <= (reset /= '1') and ( state_cur(362) or ( state_cur(361) and (NOT(in1)) = '1' ) );
	state_next(362) <= (reset /= '1') and ( ( state_cur(363) and not ( (NOT(in1)) = '1' ) ) );
	state_next(363) <= (reset /= '1') and ( state_cur(364) or ( state_cur(363) and (NOT(in1)) = '1' ) );
	state_next(364) <= (reset /= '1') and ( ( state_cur(365) and not ( (NOT(in1)) = '1' ) ) );
	state_next(365) <= (reset /= '1') and ( state_cur(366) or ( state_cur(365) and (NOT(in1)) = '1' ) );
	state_next(366) <= (reset /= '1') and ( ( state_cur(367) and not ( (NOT(in1)) = '1' ) ) );
	state_next(367) <= (reset /= '1') and ( state_cur(368) or ( state_cur(367) and (NOT(in1)) = '1' ) );
	state_next(368) <= (reset /= '1') and ( ( state_cur(369) and not ( (NOT(in1)) = '1' ) ) );
	state_next(369) <= (reset /= '1') and ( state_cur(370) or ( state_cur(369) and (NOT(in1)) = '1' ) );
	state_next(370) <= (reset /= '1') and ( ( state_cur(371) and not ( (NOT(in1)) = '1' ) ) );
	state_next(371) <= (reset /= '1') and ( state_cur(372) or ( state_cur(371) and (NOT(in1)) = '1' ) );
	state_next(372) <= (reset /= '1') and ( ( state_cur(373) and not ( (NOT(in1)) = '1' ) ) );
	state_next(373) <= (reset /= '1') and ( state_cur(374) or ( state_cur(373) and (NOT(in1)) = '1' ) );
	state_next(374) <= (reset /= '1') and ( ( state_cur(375) and not ( (NOT(in1)) = '1' ) ) );
	state_next(375) <= (reset /= '1') and ( state_cur(376) or ( state_cur(375) and (NOT(in1)) = '1' ) );
	state_next(376) <= (reset /= '1') and ( ( state_cur(377) and not ( (NOT(in1)) = '1' ) ) );
	state_next(377) <= (reset /= '1') and ( state_cur(378) or ( state_cur(377) and (NOT(in1)) = '1' ) );
	state_next(378) <= (reset /= '1') and ( ( state_cur(379) and not ( (NOT(in1)) = '1' ) ) );
	state_next(379) <= (reset /= '1') and ( state_cur(380) or ( state_cur(379) and (NOT(in1)) = '1' ) );
	state_next(380) <= (reset /= '1') and ( ( state_cur(381) and not ( (NOT(in1)) = '1' ) ) );
	state_next(381) <= (reset /= '1') and ( state_cur(382) or ( state_cur(381) and (NOT(in1)) = '1' ) );
	state_next(382) <= (reset /= '1') and ( ( state_cur(383) and not ( (NOT(in1)) = '1' ) ) );
	state_next(383) <= (reset /= '1') and ( state_cur(384) or ( state_cur(383) and (NOT(in1)) = '1' ) );
	state_next(384) <= (reset /= '1') and ( ( state_cur(385) and not ( (NOT(in1)) = '1' ) ) );
	state_next(385) <= (reset /= '1') and ( state_cur(386) or ( state_cur(385) and (NOT(in1)) = '1' ) );
	state_next(386) <= (reset /= '1') and ( ( state_cur(387) and not ( (NOT(in1)) = '1' ) ) );
	state_next(387) <= (reset /= '1') and ( state_cur(388) or ( state_cur(387) and (NOT(in1)) = '1' ) );
	state_next(388) <= (reset /= '1') and ( ( state_cur(389) and not ( (NOT(in1)) = '1' ) ) );
	state_next(389) <= (reset /= '1') and ( state_cur(390) or ( state_cur(389) and (NOT(in1)) = '1' ) );
	state_next(390) <= (reset /= '1') and ( ( state_cur(391) and not ( (NOT(in1)) = '1' ) ) );
	state_next(391) <= (reset /= '1') and ( state_cur(392) or ( state_cur(391) and (NOT(in1)) = '1' ) );
	state_next(392) <= (reset /= '1') and ( ( state_cur(393) and not ( (NOT(in1)) = '1' ) ) );
	state_next(393) <= (reset /= '1') and ( state_cur(394) or ( state_cur(393) and (NOT(in1)) = '1' ) );
	state_next(394) <= (reset /= '1') and ( ( state_cur(395) and not ( (NOT(in1)) = '1' ) ) );
	state_next(395) <= (reset /= '1') and ( state_cur(396) or ( state_cur(395) and (NOT(in1)) = '1' ) );
	state_next(396) <= (reset /= '1') and ( ( state_cur(397) and not ( (NOT(in1)) = '1' ) ) );
	state_next(397) <= (reset /= '1') and ( state_cur(398) or ( state_cur(397) and (NOT(in1)) = '1' ) );
	state_next(398) <= (reset /= '1') and ( ( state_cur(399) and not ( (NOT(in1)) = '1' ) ) );
	state_next(399) <= (reset /= '1') and ( state_cur(400) or ( state_cur(399) and (NOT(in1)) = '1' ) );
	state_next(400) <= (reset /= '1') and ( ( state_cur(401) and not ( (NOT(in1)) = '1' ) ) );
	state_next(401) <= (reset /= '1') and ( state_cur(402) or ( state_cur(401) and (NOT(in1)) = '1' ) );
	state_next(402) <= (reset /= '1') and ( ( state_cur(403) and not ( (NOT(in1)) = '1' ) ) );
	state_next(403) <= (reset /= '1') and ( state_cur(404) or ( state_cur(403) and (NOT(in1)) = '1' ) );
	state_next(404) <= (reset /= '1') and ( ( state_cur(405) and not ( (NOT(in1)) = '1' ) ) );
	state_next(405) <= (reset /= '1') and ( state_cur(406) or ( state_cur(405) and (NOT(in1)) = '1' ) );
	state_next(406) <= (reset /= '1') and ( ( state_cur(407) and not ( (NOT(in1)) = '1' ) ) );
	state_next(407) <= (reset /= '1') and ( state_cur(408) or ( state_cur(407) and (NOT(in1)) = '1' ) );
	state_next(408) <= (reset /= '1') and ( ( state_cur(409) and not ( (NOT(in1)) = '1' ) ) );
	state_next(409) <= (reset /= '1') and ( state_cur(410) or ( state_cur(409) and (NOT(in1)) = '1' ) );
	state_next(410) <= (reset /= '1') and ( ( state_cur(411) and not ( (NOT(in1)) = '1' ) ) );
	state_next(411) <= (reset /= '1') and ( state_cur(412) or ( state_cur(411) and (NOT(in1)) = '1' ) );
	state_next(412) <= (reset /= '1') and ( ( state_cur(413) and not ( (NOT(in1)) = '1' ) ) );
	state_next(413) <= (reset /= '1') and ( state_cur(414) or ( state_cur(413) and (NOT(in1)) = '1' ) );
	state_next(414) <= (reset /= '1') and ( ( state_cur(415) and not ( (NOT(in1)) = '1' ) ) );
	state_next(415) <= (reset /= '1') and ( state_cur(416) or ( state_cur(415) and (NOT(in1)) = '1' ) );
	state_next(416) <= (reset /= '1') and ( ( state_cur(417) and not ( (NOT(in1)) = '1' ) ) );
	state_next(417) <= (reset /= '1') and ( state_cur(418) or ( state_cur(417) and (NOT(in1)) = '1' ) );
	state_next(418) <= (reset /= '1') and ( ( state_cur(419) and not ( (NOT(in1)) = '1' ) ) );
	state_next(419) <= (reset /= '1') and ( state_cur(420) or ( state_cur(419) and (NOT(in1)) = '1' ) );
	state_next(420) <= (reset /= '1') and ( ( state_cur(421) and not ( (NOT(in1)) = '1' ) ) );
	state_next(421) <= (reset /= '1') and ( state_cur(422) or ( state_cur(421) and (NOT(in1)) = '1' ) );
	state_next(422) <= (reset /= '1') and ( ( state_cur(423) and not ( (NOT(in1)) = '1' ) ) );
	state_next(423) <= (reset /= '1') and ( state_cur(424) or ( state_cur(423) and (NOT(in1)) = '1' ) );
	state_next(424) <= (reset /= '1') and ( ( state_cur(425) and not ( (NOT(in1)) = '1' ) ) );
	state_next(425) <= (reset /= '1') and ( state_cur(426) or ( state_cur(425) and (NOT(in1)) = '1' ) );
	state_next(426) <= (reset /= '1') and ( ( state_cur(427) and not ( (NOT(in1)) = '1' ) ) );
	state_next(427) <= (reset /= '1') and ( state_cur(428) or ( state_cur(427) and (NOT(in1)) = '1' ) );
	state_next(428) <= (reset /= '1') and ( ( state_cur(429) and not ( (NOT(in1)) = '1' ) ) );
	state_next(429) <= (reset /= '1') and ( state_cur(430) or ( state_cur(429) and (NOT(in1)) = '1' ) );
	state_next(430) <= (reset /= '1') and ( ( state_cur(431) and not ( (NOT(in1)) = '1' ) ) );
	state_next(431) <= (reset /= '1') and ( state_cur(432) or ( state_cur(431) and (NOT(in1)) = '1' ) );
	state_next(432) <= (reset /= '1') and ( ( state_cur(433) and not ( (NOT(in1)) = '1' ) ) );
	state_next(433) <= (reset /= '1') and ( state_cur(434) or ( state_cur(433) and (NOT(in1)) = '1' ) );
	state_next(434) <= (reset /= '1') and ( ( state_cur(435) and not ( (NOT(in1)) = '1' ) ) );
	state_next(435) <= (reset /= '1') and ( state_cur(436) or ( state_cur(435) and (NOT(in1)) = '1' ) );
	state_next(436) <= (reset /= '1') and ( ( state_cur(437) and not ( (NOT(in1)) = '1' ) ) );
	state_next(437) <= (reset /= '1') and ( state_cur(438) or ( state_cur(437) and (NOT(in1)) = '1' ) );
	state_next(438) <= (reset /= '1') and ( ( state_cur(439) and not ( (NOT(in1)) = '1' ) ) );
	state_next(439) <= (reset /= '1') and ( state_cur(440) or ( state_cur(439) and (NOT(in1)) = '1' ) );
	state_next(440) <= (reset /= '1') and ( ( state_cur(441) and not ( (NOT(in1)) = '1' ) ) );
	state_next(441) <= (reset /= '1') and ( state_cur(442) or ( state_cur(441) and (NOT(in1)) = '1' ) );
	state_next(442) <= (reset /= '1') and ( ( state_cur(443) and not ( (NOT(in1)) = '1' ) ) );
	state_next(443) <= (reset /= '1') and ( state_cur(444) or ( state_cur(443) and (NOT(in1)) = '1' ) );
	state_next(444) <= (reset /= '1') and ( ( state_cur(445) and not ( (NOT(in1)) = '1' ) ) );
	state_next(445) <= (reset /= '1') and ( state_cur(446) or ( state_cur(445) and (NOT(in1)) = '1' ) );
	state_next(446) <= (reset /= '1') and ( ( state_cur(447) and not ( (NOT(in1)) = '1' ) ) );
	state_next(447) <= (reset /= '1') and ( state_cur(448) or ( state_cur(447) and (NOT(in1)) = '1' ) );
	state_next(448) <= (reset /= '1') and ( ( state_cur(449) and not ( (NOT(in1)) = '1' ) ) );
	state_next(449) <= (reset /= '1') and ( state_cur(450) or ( state_cur(449) and (NOT(in1)) = '1' ) );
	state_next(450) <= (reset /= '1') and ( ( state_cur(451) and not ( (NOT(in1)) = '1' ) ) );
	state_next(451) <= (reset /= '1') and ( state_cur(452) or ( state_cur(451) and (NOT(in1)) = '1' ) );
	state_next(452) <= (reset /= '1') and ( ( state_cur(453) and not ( (NOT(in1)) = '1' ) ) );
	state_next(453) <= (reset /= '1') and ( state_cur(454) or ( state_cur(453) and (NOT(in1)) = '1' ) );
	state_next(454) <= (reset /= '1') and ( ( state_cur(455) and not ( (NOT(in1)) = '1' ) ) );
	state_next(455) <= (reset /= '1') and ( state_cur(456) or ( state_cur(455) and (NOT(in1)) = '1' ) );
	state_next(456) <= (reset /= '1') and ( ( state_cur(457) and not ( (NOT(in1)) = '1' ) ) );
	state_next(457) <= (reset /= '1') and ( state_cur(458) or ( state_cur(457) and (NOT(in1)) = '1' ) );
	state_next(458) <= (reset /= '1') and ( ( state_cur(459) and not ( (NOT(in1)) = '1' ) ) );
	state_next(459) <= (reset /= '1') and ( state_cur(460) or ( state_cur(459) and (NOT(in1)) = '1' ) );
	state_next(460) <= (reset /= '1') and ( ( state_cur(461) and not ( (NOT(in1)) = '1' ) ) );
	state_next(461) <= (reset /= '1') and ( state_cur(462) or ( state_cur(461) and (NOT(in1)) = '1' ) );
	state_next(462) <= (reset /= '1') and ( ( state_cur(463) and not ( (NOT(in1)) = '1' ) ) );
	state_next(463) <= (reset /= '1') and ( state_cur(464) or ( state_cur(463) and (NOT(in1)) = '1' ) );
	state_next(464) <= (reset /= '1') and ( ( state_cur(465) and not ( (NOT(in1)) = '1' ) ) );
	state_next(465) <= (reset /= '1') and ( state_cur(466) or ( state_cur(465) and (NOT(in1)) = '1' ) );
	state_next(466) <= (reset /= '1') and ( ( state_cur(467) and not ( (NOT(in1)) = '1' ) ) );
	state_next(467) <= (reset /= '1') and ( state_cur(468) or ( state_cur(467) and (NOT(in1)) = '1' ) );
	state_next(468) <= (reset /= '1') and ( ( state_cur(469) and not ( (NOT(in1)) = '1' ) ) );
	state_next(469) <= (reset /= '1') and ( state_cur(470) or ( state_cur(469) and (NOT(in1)) = '1' ) );
	state_next(470) <= (reset /= '1') and ( ( state_cur(471) and not ( (NOT(in1)) = '1' ) ) );
	state_next(471) <= (reset /= '1') and ( state_cur(472) or ( state_cur(471) and (NOT(in1)) = '1' ) );
	state_next(472) <= (reset /= '1') and ( ( state_cur(473) and not ( (NOT(in1)) = '1' ) ) );
	state_next(473) <= (reset /= '1') and ( state_cur(474) or ( state_cur(473) and (NOT(in1)) = '1' ) );
	state_next(474) <= (reset /= '1') and ( ( state_cur(475) and not ( (NOT(in1)) = '1' ) ) );
	state_next(475) <= (reset /= '1') and ( state_cur(476) or ( state_cur(475) and (NOT(in1)) = '1' ) );
	state_next(476) <= (reset /= '1') and ( ( state_cur(477) and not ( (NOT(in1)) = '1' ) ) );
	state_next(477) <= (reset /= '1') and ( state_cur(478) or ( state_cur(477) and (NOT(in1)) = '1' ) );
	state_next(478) <= (reset /= '1') and ( ( state_cur(479) and not ( (NOT(in1)) = '1' ) ) );
	state_next(479) <= (reset /= '1') and ( state_cur(480) or ( state_cur(479) and (NOT(in1)) = '1' ) );
	state_next(480) <= (reset /= '1') and ( ( state_cur(481) and not ( (NOT(in1)) = '1' ) ) );
	state_next(481) <= (reset /= '1') and ( state_cur(482) or ( state_cur(481) and (NOT(in1)) = '1' ) );
	state_next(482) <= (reset /= '1') and ( ( state_cur(483) and not ( (NOT(in1)) = '1' ) ) );
	state_next(483) <= (reset /= '1') and ( state_cur(484) or ( state_cur(483) and (NOT(in1)) = '1' ) );
	state_next(484) <= (reset /= '1') and ( ( state_cur(485) and not ( (NOT(in1)) = '1' ) ) );
	state_next(485) <= (reset /= '1') and ( state_cur(486) or ( state_cur(485) and (NOT(in1)) = '1' ) );
	state_next(486) <= (reset /= '1') and ( ( state_cur(487) and not ( (NOT(in1)) = '1' ) ) );
	state_next(487) <= (reset /= '1') and ( state_cur(488) or ( state_cur(487) and (NOT(in1)) = '1' ) );
	state_next(488) <= (reset /= '1') and ( ( state_cur(489) and not ( (NOT(in1)) = '1' ) ) );
	state_next(489) <= (reset /= '1') and ( state_cur(490) or ( state_cur(489) and (NOT(in1)) = '1' ) );
	state_next(490) <= (reset /= '1') and ( ( state_cur(491) and not ( (NOT(in1)) = '1' ) ) );
	state_next(491) <= (reset /= '1') and ( state_cur(492) or ( state_cur(491) and (NOT(in1)) = '1' ) );
	state_next(492) <= (reset /= '1') and ( ( state_cur(493) and not ( (NOT(in1)) = '1' ) ) );
	state_next(493) <= (reset /= '1') and ( state_cur(494) or ( state_cur(493) and (NOT(in1)) = '1' ) );
	state_next(494) <= (reset /= '1') and ( ( state_cur(495) and not ( (NOT(in1)) = '1' ) ) );
	state_next(495) <= (reset /= '1') and ( state_cur(496) or ( state_cur(495) and (NOT(in1)) = '1' ) );
	state_next(496) <= (reset /= '1') and ( ( state_cur(497) and not ( (NOT(in1)) = '1' ) ) );
	state_next(497) <= (reset /= '1') and ( state_cur(498) or ( state_cur(497) and (NOT(in1)) = '1' ) );
	state_next(498) <= (reset /= '1') and ( ( state_cur(499) and not ( (NOT(in1)) = '1' ) ) );
	state_next(499) <= (reset /= '1') and ( state_cur(500) or ( state_cur(499) and (NOT(in1)) = '1' ) );
	state_next(500) <= (reset /= '1') and ( ( state_cur(501) and not ( (NOT(in1)) = '1' ) ) );
	state_next(501) <= (reset /= '1') and ( state_cur(502) or ( state_cur(501) and (NOT(in1)) = '1' ) );
	state_next(502) <= (reset /= '1') and ( ( state_cur(503) and not ( (NOT(in1)) = '1' ) ) );
	state_next(503) <= (reset /= '1') and ( state_cur(504) or ( state_cur(503) and (NOT(in1)) = '1' ) );
	state_next(504) <= (reset /= '1') and ( ( state_cur(505) and not ( (NOT(in1)) = '1' ) ) );
	state_next(505) <= (reset /= '1') and ( state_cur(506) or ( state_cur(505) and (NOT(in1)) = '1' ) );
	state_next(506) <= (reset /= '1') and ( ( state_cur(507) and not ( (NOT(in1)) = '1' ) ) );
	state_next(507) <= (reset /= '1') and ( state_cur(508) or ( state_cur(507) and (NOT(in1)) = '1' ) );
	state_next(508) <= (reset /= '1') and ( ( state_cur(509) and not ( (NOT(in1)) = '1' ) ) );
	state_next(509) <= (reset /= '1') and ( state_cur(510) or ( state_cur(509) and (NOT(in1)) = '1' ) );
	state_next(510) <= (reset /= '1') and ( ( state_cur(511) and not ( (NOT(in1)) = '1' ) ) );
	state_next(511) <= (reset /= '1') and ( state_cur(512) or ( state_cur(511) and (NOT(in1)) = '1' ) );
	state_next(512) <= (reset /= '1') and ( ( state_cur(513) and not ( (NOT(in1)) = '1' ) ) );
	state_next(513) <= (reset /= '1') and ( state_cur(514) or ( state_cur(513) and (NOT(in1)) = '1' ) );
	state_next(514) <= (reset /= '1') and ( ( state_cur(515) and not ( (NOT(in1)) = '1' ) ) );
	state_next(515) <= (reset /= '1') and ( state_cur(516) or ( state_cur(515) and (NOT(in1)) = '1' ) );
	state_next(516) <= (reset /= '1') and ( ( state_cur(517) and not ( (NOT(in1)) = '1' ) ) );
	state_next(517) <= (reset /= '1') and ( state_cur(518) or ( state_cur(517) and (NOT(in1)) = '1' ) );
	state_next(518) <= (reset /= '1') and ( ( state_cur(519) and not ( (NOT(in1)) = '1' ) ) );
	state_next(519) <= (reset /= '1') and ( ( state_cur(519) and (NOT(in1)) = '1' ) or state_cur(1) );
	state_next(520) <= (reset /= '1') and ( ( state_cur(520) and (NOT(in1)) = '1' ) or state_cur(73) );
	state_next(521) <= (reset /= '1') and ( ( state_cur(521) and (NOT(in1)) = '1' ) or state_cur(71) );
	state_next(522) <= (reset /= '1') and ( ( state_cur(220) and not ( (in6) = '1' ) ) );
	state_next(523) <= (reset /= '1') and ( state_cur(149) );

	-- Assignment of buffers for buffered outputs

	out386_bufn <= state_cur(186) or state_cur(270);
	out404_bufn <= (state_cur(290) = '1' and rtmcmp290 = '0') or state_cur(291) or state_cur(173);
	out457_bufn <= state_cur(142) or state_cur(190) or state_cur(169);
	out841_bufn <= rtmcmp92 or state_cur(189);
	out276_bufn <= state_cur(233) or state_cur(274);
	out67_bufn <= state_cur(189) or state_cur(282) or state_cur(98) or state_cur(203) or (state_cur(92) = '1' and rtmcmp92 = '0') or state_cur(336) or state_cur(337);
	out239_bufn <= ( state_cur(240) and (in7) = '1' ) or state_cur(523) or state_cur(129);
	out259_bufn <= state_cur(268) or state_cur(178) or ( state_cur(220) and (in6) = '1' ) or ( state_cur(150) and (in3) = '1' ) or ( state_cur(175) and (in4) = '1' ) or ( state_cur(208) and (in5) = '1' ) or state_cur(523) or state_cur(129);
	out416_bufn <= state_cur(338) or state_cur(143) or state_cur(289) or state_cur(322);
	out646_bufn <= state_cur(340) or state_cur(326);
	out485_bufn <= ( state_cur(240) and (in7) = '1' ) or ( state_cur(150) and (in3) = '1' );
	out935_bufn <= state_cur(193) or state_cur(134);
	out463_bufn <= state_cur(338) or state_cur(119) or state_cur(134) or state_cur(233) or state_cur(174);
	out120_bufn <= rtmcmp92 or state_cur(100) or state_cur(91) or state_cur(179) or state_cur(228);
	out293_bufn <= state_cur(342) or state_cur(303);
	out216_bufn <= state_cur(107) or state_cur(212) or rtmcmp128 or (state_cur(276) = '1' and rtmcmp276 = '0') or state_cur(114) or state_cur(326) or state_cur(123) or state_cur(190) or state_cur(186) or rtmcmp290 or state_cur(204) or state_cur(191) or state_cur(303) or rtmcmp276;
	out319_bufn <= (state_cur(276) = '1' and rtmcmp276 = '0') or state_cur(114) or state_cur(99) or state_cur(218) or (state_cur(128) = '1' and rtmcmp128 = '0') or state_cur(296);
	out230_bufn <= ( state_cur(220) and (in6) = '1' ) or state_cur(224);
	out1_bufn <= ( state_cur(317) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(305) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(215) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(316) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(121) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(84) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(122) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(192) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(194) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(295) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(313) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(264) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(10) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(67) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(75) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(28) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(243) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(87) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(124) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(240) and not ( (in7) = '1' ) ) or ( state_cur(269) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(50) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(64) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(68) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(49) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(171) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(130) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(77) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(302) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(287) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(176) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(216) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(250) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(202) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(318) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(136) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(211) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(120) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(135) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(226) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(279) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(55) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(167) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(165) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(163) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(161) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(159) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(157) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(155) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(101) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(116) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(118) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(127) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(314) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(304) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(112) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(140) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(288) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(217) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(80) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(272) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(297) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(278) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(258) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(256) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(24) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(65) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(246) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(61) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(12) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(104) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(21) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(51) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(52) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(46) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(37) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(41) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(285) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(323) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(35) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(34) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(259) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(33) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(324) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(320) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(117) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(26) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(27) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(14) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(239) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(188) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(263) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(13) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(17) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(207) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(6) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(48) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(201) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(44) and not ( (NOT(in0)) = '1' ) ) or ( state_cur(90) and not ( (NOT(in0)) = '1' ) );
	out93_bufn <= state_cur(522) or state_cur(93) or state_cur(96) or state_cur(108) or ( state_cur(220) and (in6) = '1' ) or state_cur(342) or state_cur(340) or state_cur(95) or state_cur(184) or ( state_cur(150) and (in3) = '1' ) or state_cur(187) or ( state_cur(175) and (in4) = '1' ) or ( state_cur(208) and (in5) = '1' ) or state_cur(334) or state_cur(339);
	out89_bufn <= state_cur(149) or state_cur(341) or state_cur(522) or state_cur(93) or state_cur(94) or state_cur(96) or state_cur(213) or state_cur(108) or state_cur(281) or state_cur(103) or state_cur(342) or state_cur(340) or state_cur(95) or state_cur(184) or state_cur(183) or state_cur(280) or state_cur(187) or state_cur(331) or state_cur(224) or state_cur(301) or state_cur(200) or state_cur(333) or state_cur(334) or state_cur(339);
	out539_bufn <= state_cur(142) or state_cur(190);
	out62_bufn <= state_cur(193) or rtmcmp92 or state_cur(107) or state_cur(212) or state_cur(338) or state_cur(119) or rtmcmp128 or state_cur(100) or (state_cur(276) = '1' and rtmcmp276 = '0') or state_cur(114) or state_cur(134) or state_cur(236) or state_cur(189) or state_cur(326) or state_cur(312) or state_cur(123) or state_cur(91) or state_cur(233) or state_cur(190) or state_cur(186) or state_cur(179) or rtmcmp290 or state_cur(282) or state_cur(319) or state_cur(174) or state_cur(204) or state_cur(172) or state_cur(191) or state_cur(303) or state_cur(274) or rtmcmp276 or state_cur(98) or state_cur(203) or state_cur(228) or (state_cur(92) = '1' and rtmcmp92 = '0') or state_cur(336) or state_cur(337);
	out856_bufn <= state_cur(107) or state_cur(147) or state_cur(236);
	out451_bufn <= state_cur(123) or state_cur(169);
	out287_bufn <= state_cur(332) or state_cur(303);
	out315_bufn <= state_cur(268) or state_cur(178) or (state_cur(128) = '1' and rtmcmp128 = '0') or state_cur(296);
	out536_bufn <= state_cur(95) or state_cur(190);
	out209_bufn <= state_cur(191) or state_cur(200);
	out221_bufn <= rtmcmp128 or state_cur(237) or state_cur(197) or rtmcmp276;
	out283_bufn <= state_cur(193) or state_cur(236) or state_cur(312) or state_cur(319) or state_cur(172) or state_cur(274);
	out368_bufn <= state_cur(213) or ( state_cur(175) and (in4) = '1' );
	out516_bufn <= ( state_cur(208) and not ( (in5) = '1' ) ) or state_cur(281) or state_cur(183) or state_cur(280);
	out393_bufn <= state_cur(193) or state_cur(212) or state_cur(338) or state_cur(143) or state_cur(210) or state_cur(289) or state_cur(322) or state_cur(204);
	out1008_bufn <= state_cur(182) or state_cur(268) or state_cur(178);
	out392_bufn <= state_cur(108) or state_cur(204);
	out261_bufn <= state_cur(268) or state_cur(178) or state_cur(523) or state_cur(129);
	out559_bufn <= state_cur(99) or state_cur(218);
	out543_bufn <= state_cur(326) or state_cur(292) or state_cur(123) or state_cur(233);
	out895_bufn <= state_cur(219) or state_cur(125) or state_cur(247) or state_cur(242) or state_cur(241) or state_cur(148);
	out82_bufn <= ( state_cur(208) and (in5) = '1' ) or (state_cur(92) = '1' and rtmcmp92 = '0') or state_cur(336);
	out220_bufn <= state_cur(107) or rtmcmp128 or state_cur(147) or state_cur(237) or state_cur(236) or state_cur(197) or rtmcmp276;
	out95_bufn <= state_cur(522) or state_cur(93) or state_cur(96) or state_cur(108) or state_cur(342) or state_cur(340) or state_cur(95) or state_cur(184) or state_cur(187) or state_cur(334) or state_cur(339);
	out943_bufn <= (state_cur(290) = '1' and rtmcmp290 = '0') or state_cur(291) or (state_cur(276) = '1' and rtmcmp276 = '0') or state_cur(114);
	out465_bufn <= state_cur(319) or state_cur(174);
	out238_bufn <= ( state_cur(175) and (in4) = '1' ) or state_cur(523) or state_cur(129);
	out1025_bufn <= ( state_cur(328) and (in11) = '1' ) or state_cur(268) or state_cur(178);
	out132_bufn <= state_cur(146) or state_cur(138) or state_cur(273) or state_cur(105);
	out79_bufn <= ( state_cur(328) and (in11) = '1' ) or state_cur(98) or state_cur(228) or (state_cur(92) = '1' and rtmcmp92 = '0') or state_cur(336);
	out500_bufn <= state_cur(91) or state_cur(282);
	out65_bufn <= state_cur(179) or state_cur(337);
	out111_bufn <= state_cur(96) or state_cur(95) or state_cur(334);
	out420_bufn <= ( state_cur(328) and (in11) = '1' ) or state_cur(306);
	out1076_bufn <= state_cur(93) or state_cur(107);
	out101_bufn <= state_cur(523) or state_cur(129) or ( state_cur(175) and not ( (in4) = '1' ) );
	out106_bufn <= ( state_cur(220) and not ( (in6) = '1' ) ) or state_cur(341) or state_cur(94) or ( state_cur(150) and not ( (in3) = '1' ) ) or state_cur(213) or ( state_cur(208) and not ( (in5) = '1' ) ) or state_cur(281) or state_cur(183) or state_cur(280) or state_cur(224) or state_cur(200) or state_cur(333) or ( state_cur(175) and not ( (in4) = '1' ) );
	out68_bufn <= state_cur(193) or rtmcmp92 or state_cur(338) or state_cur(119) or state_cur(100) or state_cur(134) or state_cur(236) or state_cur(189) or state_cur(312) or state_cur(91) or state_cur(233) or state_cur(179) or state_cur(282) or state_cur(319) or state_cur(174) or state_cur(172) or state_cur(274) or state_cur(98) or state_cur(203) or state_cur(228) or (state_cur(92) = '1' and rtmcmp92 = '0') or state_cur(336) or state_cur(337);
	out1069_bufn <= state_cur(213) or state_cur(212);
	out77_bufn <= state_cur(228) or (state_cur(92) = '1' and rtmcmp92 = '0') or state_cur(336);
	out102_bufn <= state_cur(94) or state_cur(213) or ( state_cur(175) and not ( (in4) = '1' ) );
	out394_bufn <= state_cur(193) or state_cur(212) or state_cur(210) or state_cur(204);
	out342_bufn <= ( state_cur(220) and (in6) = '1' ) or ( state_cur(150) and (in3) = '1' ) or ( state_cur(175) and (in4) = '1' ) or ( state_cur(208) and (in5) = '1' );
	out104_bufn <= ( state_cur(220) and not ( (in6) = '1' ) ) or state_cur(341) or state_cur(94) or ( state_cur(150) and not ( (in3) = '1' ) ) or state_cur(213) or ( state_cur(208) and not ( (in5) = '1' ) ) or state_cur(281) or ( state_cur(220) and (in6) = '1' ) or state_cur(146) or state_cur(138) or state_cur(183) or state_cur(280) or ( state_cur(150) and (in3) = '1' ) or ( state_cur(175) and (in4) = '1' ) or ( state_cur(208) and (in5) = '1' ) or state_cur(224) or state_cur(200) or state_cur(273) or state_cur(105) or state_cur(333) or ( state_cur(175) and not ( (in4) = '1' ) );
	out361_bufn <= state_cur(338) or state_cur(172);
	out116_bufn <= ( state_cur(150) and not ( (in3) = '1' ) ) or state_cur(200) or state_cur(333);
	out595_bufn <= state_cur(119) or state_cur(237) or state_cur(236) or state_cur(312);
	out1004_bufn <= state_cur(143) or state_cur(132);
	out227_bufn <= state_cur(123) or state_cur(224);
	out109_bufn <= state_cur(186) or state_cur(334);
	out619_bufn <= state_cur(237) or state_cur(312);
	out410_bufn <= state_cur(335) or state_cur(143) or state_cur(132) or state_cur(322);
	out989_bufn <= ( state_cur(150) and not ( (in3) = '1' ) ) or ( state_cur(240) and (in7) = '1' );
	out431_bufn <= state_cur(184) or state_cur(187);
	out938_bufn <= state_cur(94) or (state_cur(276) = '1' and rtmcmp276 = '0') or state_cur(114);
	out525_bufn <= state_cur(96) or rtmcmp290;
	out73_bufn <= rtmcmp92 or (state_cur(290) = '1' and rtmcmp290 = '0') or state_cur(291) or state_cur(91) or state_cur(203) or (state_cur(92) = '1' and rtmcmp92 = '0') or state_cur(336) or state_cur(337);
	out837_bufn <= state_cur(522) or state_cur(108) or state_cur(342);
	out860_bufn <= state_cur(119) or state_cur(236);
	out228_bufn <= ( state_cur(220) and not ( (in6) = '1' ) ) or state_cur(341) or state_cur(224);
	out421_bufn <= ( state_cur(328) and (in11) = '1' ) or ( state_cur(325) and not ( (in10) = '1' ) ) or ( state_cur(97) and not ( (NOT(in0)) = '1' ) ) or state_cur(306);
	out409_bufn <= state_cur(132) or state_cur(322);
	out473_bufn <= state_cur(99) or state_cur(218) or ( state_cur(325) and (in10) = '1' ) or ( state_cur(310) and not ( (in9) = '1' ) );
	out509_bufn <= state_cur(123) or state_cur(223);
	out94_bufn <= rtmcmp276 or state_cur(339);
	out1048_bufn <= state_cur(341) or rtmcmp128;
	out98_bufn <= state_cur(93) or state_cur(340) or state_cur(339);
	out945_bufn <= ( state_cur(240) and (in7) = '1' ) or (state_cur(276) = '1' and rtmcmp276 = '0') or state_cur(114);
	out156_bufn <= ( state_cur(328) and (in11) = '1' ) or state_cur(98);
	out152_bufn <= state_cur(100) or state_cur(203);

	-- Assignment of non-buffered outputs

	out80 <=
		state_cur(92);
	out576 <=
		state_cur(200);
	out1103 <=
		state_cur(336);
	out438 <=
		state_cur(151);
	out171 <=
		state_cur(222) or state_cur(102);
	out378 <=
		state_cur(340) or state_cur(222) or state_cur(138);
	out940 <=
		state_cur(276);
	out131 <=
		state_cur(99);
	out376 <=
		state_cur(138);
	out891 <=
		state_cur(237);
	out611 <=
		state_cur(209);
	out638 <=
		state_cur(222) or state_cur(209);
	out354 <=
		state_cur(129);
	out7 <=
		state_cur(3);
	out1127 <=
		state_cur(339);
	out888 <=
		state_cur(237);
	out1141 <=
		state_cur(348);
	out6 <=
		state_cur(2);
	out1200 <=
		state_cur(466);
	out1148 <=
		state_cur(362);
	out250 <=
		state_cur(114);
	out1100 <=
		state_cur(335);
	out1168 <=
		state_cur(402);
	out1158 <=
		state_cur(382);
	out581 <=
		state_cur(204);
	out549 <=
		state_cur(222) or state_cur(193);
	out412 <=
		state_cur(145);
	out381 <=
		state_cur(222) or state_cur(213) or state_cur(138);
	out38 <=
		state_cur(56);
	out100 <=
		state_cur(522) or state_cur(342) or state_cur(341) or state_cur(340) or state_cur(339) or state_cur(334) or state_cur(333) or state_cur(331) or
		state_cur(301) or state_cur(281) or state_cur(280) or state_cur(224) or state_cur(213) or state_cur(200) or state_cur(187) or state_cur(184) or
		state_cur(183) or state_cur(149) or state_cur(108) or state_cur(103) or state_cur(96) or state_cur(95) or state_cur(94) or state_cur(93);
	out1181 <=
		state_cur(428);
	out22 <=
		state_cur(20);
	out56 <=
		state_cur(85);
	out224 <=
		state_cur(326) or state_cur(303) or state_cur(292) or rtmcmp276 or state_cur(237) or state_cur(236) or state_cur(233) or state_cur(197) or
		state_cur(147) or rtmcmp128 or state_cur(123) or state_cur(107);
	out1115 <=
		state_cur(336);
	out191 <=
		state_cur(102);
	out290 <=
		state_cur(123);
	out1226 <=
		state_cur(518);
	out921 <=
		state_cur(271);
	out535 <=
		state_cur(191);
	out489 <=
		state_cur(178);
	out13 <=
		state_cur(8);
	out1161 <=
		state_cur(388);
	out408 <=
		state_cur(144);
	out1197 <=
		state_cur(460);
	out521 <=
		state_cur(184);
	out128 <=
		state_cur(296) or state_cur(218) or state_cur(114) or state_cur(99);
	out440 <=
		state_cur(154);
	out330 <=
		state_cur(128);
	out1003 <=
		state_cur(294);
	out1145 <=
		state_cur(356);
	out1156 <=
		state_cur(378);
	out497 <=
		state_cur(268) or state_cur(222) or state_cur(178);
	out52 <=
		state_cur(79);
	out659 <=
		state_cur(218);
	out566 <=
		state_cur(197);
	out850 <=
		state_cur(231);
	out1123 <=
		state_cur(338);
	out558 <=
		state_cur(197);
	out902 <=
		state_cur(248);
	out1217 <=
		state_cur(500);
	out357 <=
		state_cur(132);
	out229 <=
		state_cur(108);
	out1096 <=
		state_cur(335);
	out1188 <=
		state_cur(442);
	out39 <=
		state_cur(57);
	out118 <=
		state_cur(96);
	out387 <=
		state_cur(142);
	out514 <=
		state_cur(183);
	out425 <=
		state_cur(148);
	out508 <=
		state_cur(182);
	out1155 <=
		state_cur(376);
	out877 <=
		state_cur(236);
	out844 <=
		state_cur(228);
	out237 <=
		state_cur(113);
	out1133 <=
		state_cur(341);
	out1046 <=
		state_cur(301);
	out365 <=
		state_cur(137);
	out858 <=
		state_cur(233);
	out873 <=
		state_cur(235);
	out909 <=
		state_cur(260);
	out846 <=
		state_cur(230);
	out484 <=
		state_cur(177);
	out836 <=
		state_cur(224);
	out898 <=
		state_cur(242);
	out1196 <=
		state_cur(458);
	out26 <=
		state_cur(30);
	out1147 <=
		state_cur(360);
	out744 <=
		state_cur(342) or state_cur(273) or state_cur(222);
	out1026 <=
		state_cur(296);
	out430 <=
		state_cur(149);
	out962 <=
		state_cur(281);
	out45 <=
		state_cur(66);
	out9 <=
		state_cur(5);
	out1002 <=
		state_cur(294);
	out1139 <=
		state_cur(344);
	out1143 <=
		state_cur(352);
	out1173 <=
		state_cur(412);
	out28 <=
		state_cur(32);
	out1092 <=
		state_cur(334);
	out1140 <=
		state_cur(346);
	out40 <=
		state_cur(58);
	out119 <=
		state_cur(98);
	out382 <=
		state_cur(139);
	out241 <=
		state_cur(114);
	out91 <=
		state_cur(93);
	out920 <=
		state_cur(270);
	out986 <=
		state_cur(290);
	out657 <=
		state_cur(222) or state_cur(218);
	out375 <=
		state_cur(331) or state_cur(222) or state_cur(138);
	out866 <=
		state_cur(235);
	out577 <=
		state_cur(203);
	out1159 <=
		state_cur(384);
	out236 <=
		state_cur(111);
	out367 <=
		state_cur(339) or state_cur(222) or state_cur(138);
	out1130 <=
		state_cur(340);
	out25 <=
		state_cur(25);
	out258 <=
		state_cur(222) or state_cur(114);
	out990 <=
		state_cur(291);
	out900 <=
		state_cur(244);
	out748 <=
		state_cur(273) or state_cur(224) or state_cur(222);
	out1219 <=
		state_cur(504);
	out552 <=
		state_cur(196);
	out852 <=
		state_cur(232);
	out644 <=
		state_cur(222) or state_cur(210);
	out4 <=
		state_cur(1);
	out1142 <=
		state_cur(350);
	out1089 <=
		state_cur(333);
	out937 <=
		state_cur(275);
	out291 <=
		state_cur(335) or state_cur(332) or state_cur(303) or state_cur(169) or rtmcmp128 or state_cur(123);
	out482 <=
		state_cur(222) or state_cur(175);
	out924 <=
		state_cur(273);
	out1218 <=
		state_cur(502);
	out590 <=
		state_cur(205);
	out20 <=
		state_cur(18);
	out114 <=
		state_cur(222) or state_cur(178) or state_cur(96);
	out30 <=
		state_cur(38);
	out1224 <=
		state_cur(514);
	out107 <=
		state_cur(95);
	out915 <=
		state_cur(268);
	out34 <=
		state_cur(45);
	out1213 <=
		state_cur(492);
	out33 <=
		state_cur(43);
	out530 <=
		state_cur(187);
	out1191 <=
		state_cur(448);
	out223 <=
		state_cur(107);
	out834 <=
		state_cur(231) or state_cur(223);
	out1038 <=
		state_cur(298);
	out454 <=
		state_cur(170);
	out1087 <=
		state_cur(332);
	out233 <=
		state_cur(109);
	out66 <=
		state_cur(91);
	out347 <=
		state_cur(222) or state_cur(149) or state_cur(129);
	out848 <=
		state_cur(231);
	out746 <=
		state_cur(301) or state_cur(273) or state_cur(222);
	out695 <=
		state_cur(232) or state_cur(222);
	out1203 <=
		state_cur(472);
	out1085 <=
		state_cur(332);
	out1157 <=
		state_cur(380);
	out1039 <=
		state_cur(298);
	out532 <=
		state_cur(189);
	out1138 <=
		state_cur(342);
	out441 <=
		state_cur(156);
	out845 <=
		state_cur(229);
	out48 <=
		state_cur(71);
	out593 <=
		state_cur(222) or state_cur(208);
	out1182 <=
		state_cur(430);
	out57 <=
		state_cur(88);
	out44 <=
		state_cur(63);
	out1183 <=
		state_cur(432);
	out29 <=
		state_cur(36);
	out1015 <=
		state_cur(296);
	out910 <=
		state_cur(261);
	out524 <=
		state_cur(186);
	out958 <=
		state_cur(280);
	out460 <=
		state_cur(300) or state_cur(204) or state_cur(191) or state_cur(170);
	out50 <=
		state_cur(74);
	out304 <=
		state_cur(126);
	out130 <=
		state_cur(222) or state_cur(99);
	out833 <=
		state_cur(223);
	out513 <=
		rtmcmp290 or state_cur(223) or state_cur(182);
	out1210 <=
		state_cur(486);
	out370 <=
		state_cur(222) or state_cur(146) or state_cur(138);
	out481 <=
		state_cur(175);
	out207 <=
		state_cur(103);
	out445 <=
		state_cur(164);
	out362 <=
		state_cur(134);
	out908 <=
		state_cur(257);
	out1186 <=
		state_cur(438);
	out466 <=
		state_cur(172);
	out1083 <=
		state_cur(331);
	out475 <=
		state_cur(173);
	out19 <=
		state_cur(16);
	out645 <=
		state_cur(212);
	out582 <=
		state_cur(222) or state_cur(204);
	out547 <=
		state_cur(193);
	out1154 <=
		state_cur(374);
	out854 <=
		state_cur(232);
	out208 <=
		state_cur(222) or state_cur(178) or state_cur(103);
	out975 <=
		state_cur(286);
	out1150 <=
		state_cur(366);
	out503 <=
		state_cur(179);
	out650 <=
		state_cur(213);
	out863 <=
		state_cur(234);
	out1211 <=
		state_cur(488);
	out1228 <=
		state_cur(522);
	out5 <=
		state_cur(518) or state_cur(516) or state_cur(514) or state_cur(512) or state_cur(510) or state_cur(508) or state_cur(506) or state_cur(504) or
		state_cur(502) or state_cur(500) or state_cur(498) or state_cur(496) or state_cur(494) or state_cur(492) or state_cur(490) or state_cur(488) or
		state_cur(486) or state_cur(484) or state_cur(482) or state_cur(480) or state_cur(478) or state_cur(476) or state_cur(474) or state_cur(472) or
		state_cur(470) or state_cur(468) or state_cur(466) or state_cur(464) or state_cur(462) or state_cur(460) or state_cur(458) or state_cur(456) or
		state_cur(454) or state_cur(452) or state_cur(450) or state_cur(448) or state_cur(446) or state_cur(444) or state_cur(442) or state_cur(440) or
		state_cur(438) or state_cur(436) or state_cur(434) or state_cur(432) or state_cur(430) or state_cur(428) or state_cur(426) or state_cur(424) or
		state_cur(422) or state_cur(420) or state_cur(418) or state_cur(416) or state_cur(414) or state_cur(412) or state_cur(410) or state_cur(408) or
		state_cur(406) or state_cur(404) or state_cur(402) or state_cur(400) or state_cur(398) or state_cur(396) or state_cur(394) or state_cur(392) or
		state_cur(390) or state_cur(388) or state_cur(386) or state_cur(384) or state_cur(382) or state_cur(380) or state_cur(378) or state_cur(376) or
		state_cur(374) or state_cur(372) or state_cur(370) or state_cur(368) or state_cur(366) or state_cur(364) or state_cur(362) or state_cur(360) or
		state_cur(358) or state_cur(356) or state_cur(354) or state_cur(352) or state_cur(350) or state_cur(348) or state_cur(346) or state_cur(344) or
		state_cur(214) or state_cur(198) or state_cur(195) or state_cur(180) or state_cur(125) or state_cur(115) or state_cur(85) or state_cur(83) or
		state_cur(79) or state_cur(73) or state_cur(71) or state_cur(1);
	out1081 <=
		state_cur(330);
	out980 <=
		rtmcmp290;
	out533 <=
		state_cur(190);
	out338 <=
		state_cur(280) or state_cur(222) or state_cur(129);
	out32 <=
		state_cur(40);
	out1080 <=
		state_cur(329);
	out27 <=
		state_cur(31);
	out893 <=
		state_cur(238);
	out397 <=
		state_cur(143);
	out1000 <=
		state_cur(293);
	out55 <=
		state_cur(83);
	out235 <=
		state_cur(109);
	out1198 <=
		state_cur(462);
	out12 <=
		state_cur(7);
	out1221 <=
		state_cur(508);
	out277 <=
		state_cur(119);
	out1205 <=
		state_cur(476);
	out321 <=
		state_cur(338) or state_cur(322) or state_cur(319) or state_cur(298) or state_cur(289) or rtmcmp276 or state_cur(237) or state_cur(197) or
		state_cur(151) or state_cur(145) or state_cur(143) or rtmcmp128;
	out1216 <=
		state_cur(498);
	out999 <=
		state_cur(292);
	out1190 <=
		state_cur(446);
	out1078 <=
		state_cur(327);
	out17 <=
		state_cur(521) or state_cur(520) or state_cur(519) or state_cur(517) or state_cur(515) or state_cur(513) or state_cur(511) or state_cur(509) or
		state_cur(507) or state_cur(505) or state_cur(503) or state_cur(501) or state_cur(499) or state_cur(497) or state_cur(495) or state_cur(493) or
		state_cur(491) or state_cur(489) or state_cur(487) or state_cur(485) or state_cur(483) or state_cur(481) or state_cur(479) or state_cur(477) or
		state_cur(475) or state_cur(473) or state_cur(471) or state_cur(469) or state_cur(467) or state_cur(465) or state_cur(463) or state_cur(461) or
		state_cur(459) or state_cur(457) or state_cur(455) or state_cur(453) or state_cur(451) or state_cur(449) or state_cur(447) or state_cur(445) or
		state_cur(443) or state_cur(441) or state_cur(439) or state_cur(437) or state_cur(435) or state_cur(433) or state_cur(431) or state_cur(429) or
		state_cur(427) or state_cur(425) or state_cur(423) or state_cur(421) or state_cur(419) or state_cur(417) or state_cur(415) or state_cur(413) or
		state_cur(411) or state_cur(409) or state_cur(407) or state_cur(405) or state_cur(403) or state_cur(401) or state_cur(399) or state_cur(397) or
		state_cur(395) or state_cur(393) or state_cur(391) or state_cur(389) or state_cur(387) or state_cur(385) or state_cur(383) or state_cur(381) or
		state_cur(379) or state_cur(377) or state_cur(375) or state_cur(373) or state_cur(371) or state_cur(369) or state_cur(367) or state_cur(365) or
		state_cur(363) or state_cur(361) or state_cur(359) or state_cur(357) or state_cur(355) or state_cur(353) or state_cur(351) or state_cur(349) or
		state_cur(347) or state_cur(345) or state_cur(343) or state_cur(255) or state_cur(110) or state_cur(106) or state_cur(86) or state_cur(78) or
		state_cur(72) or state_cur(42) or state_cur(29) or state_cur(11);
	out1209 <=
		state_cur(484);
	out70 <=
		state_cur(337) or state_cur(336) or state_cur(282) or state_cur(228) or state_cur(203) or state_cur(189) or state_cur(179) or state_cur(102) or
		state_cur(100) or state_cur(98) or rtmcmp92 or state_cur(91);
	out1077 <=
		state_cur(326);
	out1215 <=
		state_cur(496);
	out285 <=
		state_cur(338) or state_cur(319) or state_cur(312) or state_cur(274) or state_cur(236) or state_cur(233) or state_cur(209) or state_cur(193) or
		state_cur(174) or state_cur(172) or state_cur(134) or state_cur(119);
	out1206 <=
		state_cur(478);
	out1175 <=
		state_cur(416);
	out1222 <=
		state_cur(510);
	out443 <=
		state_cur(160);
	out212 <=
		state_cur(105);
	out270 <=
		state_cur(296) or state_cur(114);
	out865 <=
		state_cur(234);
	out648 <=
		state_cur(222) or state_cur(212);
	out1176 <=
		state_cur(418);
	out1174 <=
		state_cur(414);
	out54 <=
		state_cur(82);
	out706 <=
		state_cur(296) or state_cur(222);
	out913 <=
		state_cur(266);
	out24 <=
		state_cur(23);
	out1164 <=
		state_cur(394);
	out729 <=
		state_cur(341) or state_cur(273) or state_cur(222);
	out1204 <=
		state_cur(474);
	out573 <=
		state_cur(199);
	out480 <=
		state_cur(222) or state_cur(174);
	out14 <=
		state_cur(9);
	out1073 <=
		state_cur(325);
	out974 <=
		state_cur(284);
	out358 <=
		state_cur(222) or state_cur(132);
	out504 <=
		state_cur(180);
	out21 <=
		state_cur(19);
	out37 <=
		state_cur(54);
	out541 <=
		state_cur(222) or state_cur(191);
	out1071 <=
		state_cur(322);
	out23 <=
		state_cur(22);
	out1122 <=
		state_cur(337);
	out8 <=
		state_cur(4);
	out839 <=
		state_cur(225);
	out35 <=
		state_cur(47);
	out988 <=
		state_cur(291);
	out419 <=
		state_cur(147);
	out976 <=
		state_cur(289);
	out973 <=
		state_cur(283);
	out58 <=
		state_cur(89);
	out424 <=
		state_cur(306) or state_cur(148);
	out450 <=
		state_cur(222) or state_cur(170);
	out1068 <=
		state_cur(321);
	out1170 <=
		state_cur(406);
	out1067 <=
		state_cur(319);
	out1225 <=
		state_cur(516);
	out1187 <=
		state_cur(440);
	out563 <=
		state_cur(222) or state_cur(197);
	out1178 <=
		state_cur(422);
	out31 <=
		state_cur(39);
	out51 <=
		state_cur(76);
	out1171 <=
		state_cur(408);
	out41 <=
		state_cur(59);
	out360 <=
		state_cur(133);
	out1162 <=
		state_cur(390);
	out403 <=
		state_cur(144);
	out1179 <=
		state_cur(424);
	out1212 <=
		state_cur(490);
	out1189 <=
		state_cur(444);
	out1166 <=
		state_cur(398);
	out42 <=
		state_cur(60);
	out1220 <=
		state_cur(506);
	out137 <=
		state_cur(99);
	out643 <=
		state_cur(210);
	out692 <=
		rtmcmp276 or state_cur(222);
	out43 <=
		state_cur(62);
	out972 <=
		state_cur(282);
	out472 <=
		state_cur(173);
	out505 <=
		state_cur(181);
	out934 <=
		state_cur(274);
	out1165 <=
		state_cur(396);
	out494 <=
		state_cur(334) or state_cur(222) or state_cur(178);
	out1208 <=
		state_cur(482);
	out1172 <=
		state_cur(410);
	out550 <=
		state_cur(195);
	out439 <=
		state_cur(152);
	out388 <=
		rtmcmp290 or state_cur(270) or state_cur(190) or state_cur(186) or state_cur(144) or state_cur(142);
	out1195 <=
		state_cur(456);
	out479 <=
		state_cur(174);
	out1193 <=
		state_cur(452);
	out105 <=
		state_cur(94);
	out903 <=
		state_cur(249);
	out697 <=
		state_cur(300) or state_cur(222);
	out1149 <=
		state_cur(364);
	out49 <=
		state_cur(73);
	out448 <=
		state_cur(169);
	out436 <=
		state_cur(150);
	out917 <=
		state_cur(270);
	out1064 <=
		state_cur(315);
	out912 <=
		state_cur(265);
	out592 <=
		state_cur(208);
	out1167 <=
		state_cur(400);
	out719 <=
		state_cur(237) or state_cur(222);
	out301 <=
		state_cur(125);
	out1152 <=
		state_cur(370);
	out1063 <=
		state_cur(312);
	out1230 <=
		state_cur(523);
	out46 <=
		state_cur(69);
	out47 <=
		state_cur(70);
	out351 <=
		state_cur(222) or state_cur(184) or state_cur(129);
	out1169 <=
		state_cur(404);
	out491 <=
		state_cur(222) or state_cur(200) or state_cur(178);
	out1061 <=
		state_cur(311);
	out434 <=
		state_cur(150);
	out76 <=
		state_cur(337) or state_cur(336) or state_cur(326) or state_cur(322) or state_cur(303) or state_cur(296) or state_cur(291) or rtmcmp290 or
		rtmcmp276 or state_cur(212) or state_cur(204) or state_cur(203) or state_cur(191) or state_cur(190) or state_cur(186) or state_cur(143) or
		state_cur(132) or rtmcmp128 or state_cur(123) or state_cur(114) or state_cur(107) or state_cur(100) or rtmcmp92 or state_cur(91);
	out840 <=
		state_cur(227);
	out88 <=
		state_cur(336) or state_cur(296) or state_cur(291) or rtmcmp290 or rtmcmp276 or rtmcmp128 or state_cur(114) or rtmcmp92;
	out356 <=
		state_cur(131);
	out442 <=
		state_cur(158);
	out1199 <=
		state_cur(464);
	out1043 <=
		state_cur(300);
	out11 <=
		state_cur(324) or state_cur(323) or state_cur(320) or state_cur(318) or state_cur(317) or state_cur(316) or state_cur(314) or state_cur(313) or
		state_cur(305) or state_cur(304) or state_cur(302) or state_cur(297) or state_cur(295) or state_cur(288) or state_cur(287) or state_cur(285) or
		state_cur(279) or state_cur(278) or state_cur(272) or state_cur(269) or state_cur(264) or state_cur(263) or state_cur(259) or state_cur(258) or
		state_cur(256) or state_cur(250) or state_cur(246) or state_cur(243) or state_cur(239) or state_cur(226) or state_cur(217) or state_cur(216) or
		state_cur(215) or state_cur(211) or state_cur(207) or state_cur(202) or state_cur(201) or state_cur(194) or state_cur(192) or state_cur(188) or
		state_cur(176) or state_cur(171) or state_cur(167) or state_cur(165) or state_cur(163) or state_cur(161) or state_cur(159) or state_cur(157) or
		state_cur(155) or state_cur(153) or state_cur(140) or state_cur(136) or state_cur(135) or state_cur(130) or state_cur(127) or state_cur(124) or
		state_cur(122) or state_cur(121) or state_cur(120) or state_cur(118) or state_cur(117) or state_cur(116) or state_cur(112) or state_cur(104) or
		state_cur(101) or state_cur(97) or state_cur(90) or state_cur(87) or state_cur(84) or state_cur(80) or state_cur(77) or state_cur(75) or
		state_cur(68) or state_cur(67) or state_cur(65) or state_cur(64) or state_cur(61) or state_cur(55) or state_cur(52) or state_cur(51) or
		state_cur(50) or state_cur(49) or state_cur(48) or state_cur(46) or state_cur(44) or state_cur(41) or state_cur(37) or state_cur(35) or
		state_cur(34) or state_cur(33) or state_cur(28) or state_cur(27) or state_cur(26) or state_cur(24) or state_cur(21) or state_cur(17) or
		state_cur(14) or state_cur(13) or state_cur(12) or state_cur(10) or state_cur(6);
	out591 <=
		state_cur(206);
	out1180 <=
		state_cur(426);
	out476 <=
		state_cur(291) or state_cur(173);
	out1059 <=
		state_cur(310);
	out92 <=
		state_cur(222) or state_cur(138) or state_cur(93);
	out418 <=
		state_cur(146);
	out1042 <=
		state_cur(299);
	out1057 <=
		state_cur(309);
	out213 <=
		state_cur(273) or state_cur(222) or state_cur(105);
	out444 <=
		state_cur(162);
	out1153 <=
		state_cur(372);
	out1056 <=
		state_cur(336) or state_cur(308);
	out957 <=
		state_cur(277);
	out344 <=
		state_cur(222) or state_cur(183) or state_cur(129);
	out545 <=
		state_cur(212) or state_cur(210) or state_cur(204) or state_cur(193);
	out1055 <=
		state_cur(308);
	out968 <=
		state_cur(282);
	out335 <=
		state_cur(222) or rtmcmp128;
	out226 <=
		state_cur(273) or state_cur(222) or state_cur(108);
	out905 <=
		state_cur(252);
	out1177 <=
		state_cur(420);
	out904 <=
		state_cur(251);
	out1053 <=
		state_cur(307);
	out1052 <=
		state_cur(306);
	out417 <=
		state_cur(145);
	out1201 <=
		state_cur(468);
	out1163 <=
		state_cur(392);
	out2 <=
		state_cur(330) or state_cur(329) or state_cur(327) or state_cur(321) or state_cur(315) or state_cur(311) or state_cur(309) or state_cur(307) or
		state_cur(299) or state_cur(293) or state_cur(286) or state_cur(284) or state_cur(283) or state_cur(277) or state_cur(275) or state_cur(271) or
		state_cur(267) or state_cur(266) or state_cur(265) or state_cur(262) or state_cur(261) or state_cur(260) or state_cur(257) or state_cur(254) or
		state_cur(253) or state_cur(252) or state_cur(251) or state_cur(249) or state_cur(248) or state_cur(244) or state_cur(238) or state_cur(230) or
		state_cur(229) or state_cur(227) or state_cur(225) or state_cur(221) or state_cur(206) or state_cur(205) or state_cur(199) or state_cur(185) or
		state_cur(181) or state_cur(177) or state_cur(168) or state_cur(166) or state_cur(164) or state_cur(162) or state_cur(160) or state_cur(158) or
		state_cur(156) or state_cur(154) or state_cur(139) or state_cur(137) or state_cur(133) or state_cur(131) or state_cur(126) or state_cur(113) or
		state_cur(111) or state_cur(89) or state_cur(88) or state_cur(82) or state_cur(81) or state_cur(76) or state_cur(74) or state_cur(70) or
		state_cur(69) or state_cur(66) or state_cur(63) or state_cur(62) or state_cur(60) or state_cur(59) or state_cur(58) or state_cur(57) or
		state_cur(56) or state_cur(54) or state_cur(53) or state_cur(47) or state_cur(45) or state_cur(43) or state_cur(40) or state_cur(39) or
		state_cur(38) or state_cur(36) or state_cur(32) or state_cur(31) or state_cur(30) or state_cur(25) or state_cur(23) or state_cur(22) or
		state_cur(20) or state_cur(19) or state_cur(18) or state_cur(16) or state_cur(15) or state_cur(9) or state_cur(8) or state_cur(7) or
		state_cur(5) or state_cur(4) or state_cur(3) or state_cur(2) or state_cur(0);
	out447 <=
		state_cur(168);
	out1202 <=
		state_cur(470);
	out1192 <=
		state_cur(450);
	out1050 <=
		state_cur(303);
	out1144 <=
		state_cur(354);
	out0 <=
		state_cur(0);
	out446 <=
		state_cur(166);
	out914 <=
		state_cur(267);
	out1194 <=
		state_cur(454);
	out906 <=
		state_cur(253);
	out1146 <=
		state_cur(358);
	out572 <=
		state_cur(198);
	out1223 <=
		state_cur(512);
	out53 <=
		state_cur(81);
	out36 <=
		state_cur(53);
	out355 <=
		state_cur(222) or state_cur(187) or state_cur(129);
	out1184 <=
		state_cur(434);
	out907 <=
		state_cur(254);
	out1207 <=
		state_cur(480);
	out18 <=
		state_cur(15);
	out108 <=
		state_cur(222) or state_cur(178) or state_cur(95);
	out1160 <=
		state_cur(386);
	out662 <=
		state_cur(218);
	out303 <=
		state_cur(247) or state_cur(242) or state_cur(241) or state_cur(197) or state_cur(152) or state_cur(148) or state_cur(125);
	out1214 <=
		state_cur(494);
	out1185 <=
		state_cur(436);
	out341 <=
		state_cur(523) or state_cur(222) or state_cur(129);
	out1151 <=
		state_cur(368);
	out652 <=
		state_cur(214);
	out390 <=
		state_cur(222) or state_cur(143);
	out523 <=
		state_cur(185);
	out686 <=
		state_cur(222);
	out155 <=
		state_cur(100);
	out682 <=
		state_cur(221);
	out680 <=
		state_cur(222) or state_cur(220);
	out679 <=
		state_cur(220);
	out678 <=
		state_cur(222) or state_cur(219);
	out677 <=
		state_cur(219);

	-- Assignment of buffered outputs

	out386 <= out386_buf;
	out404 <= out404_buf;
	out457 <= out457_buf;
	out841 <= out841_buf;
	out276 <= out276_buf;
	out67 <= out67_buf;
	out239 <= out239_buf;
	out259 <= out259_buf;
	out416 <= out416_buf;
	out646 <= out646_buf;
	out485 <= out485_buf;
	out935 <= out935_buf;
	out463 <= out463_buf;
	out120 <= out120_buf;
	out293 <= out293_buf;
	out216 <= out216_buf;
	out319 <= out319_buf;
	out230 <= out230_buf;
	out1 <= out1_buf;
	out93 <= out93_buf;
	out89 <= out89_buf;
	out539 <= out539_buf;
	out62 <= out62_buf;
	out856 <= out856_buf;
	out451 <= out451_buf;
	out287 <= out287_buf;
	out315 <= out315_buf;
	out536 <= out536_buf;
	out209 <= out209_buf;
	out221 <= out221_buf;
	out283 <= out283_buf;
	out368 <= out368_buf;
	out516 <= out516_buf;
	out393 <= out393_buf;
	out1008 <= out1008_buf;
	out392 <= out392_buf;
	out261 <= out261_buf;
	out559 <= out559_buf;
	out543 <= out543_buf;
	out895 <= out895_buf;
	out82 <= out82_buf;
	out220 <= out220_buf;
	out95 <= out95_buf;
	out943 <= out943_buf;
	out465 <= out465_buf;
	out238 <= out238_buf;
	out1025 <= out1025_buf;
	out132 <= out132_buf;
	out79 <= out79_buf;
	out500 <= out500_buf;
	out65 <= out65_buf;
	out111 <= out111_buf;
	out420 <= out420_buf;
	out1076 <= out1076_buf;
	out101 <= out101_buf;
	out106 <= out106_buf;
	out68 <= out68_buf;
	out1069 <= out1069_buf;
	out77 <= out77_buf;
	out102 <= out102_buf;
	out394 <= out394_buf;
	out342 <= out342_buf;
	out104 <= out104_buf;
	out361 <= out361_buf;
	out116 <= out116_buf;
	out595 <= out595_buf;
	out1004 <= out1004_buf;
	out227 <= out227_buf;
	out109 <= out109_buf;
	out619 <= out619_buf;
	out410 <= out410_buf;
	out989 <= out989_buf;
	out431 <= out431_buf;
	out938 <= out938_buf;
	out525 <= out525_buf;
	out73 <= out73_buf;
	out837 <= out837_buf;
	out860 <= out860_buf;
	out228 <= out228_buf;
	out421 <= out421_buf;
	out409 <= out409_buf;
	out473 <= out473_buf;
	out509 <= out509_buf;
	out94 <= out94_buf;
	out1048 <= out1048_buf;
	out98 <= out98_buf;
	out945 <= out945_buf;
	out156 <= out156_buf;
	out152 <= out152_buf;

	-- Retiming: the comparators

	rtmcmp92 <= '1' when state_cur(92) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp128 <= '1' when state_cur(128) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp276 <= '1' when state_cur(276) = '1' and rtmcounter0 = 1 else '0';
	rtmcmp290 <= '1' when state_cur(290) = '1' and rtmcounter0 = 1 else '0';

end architecture;

