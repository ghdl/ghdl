context is
context is