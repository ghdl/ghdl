entity tb is
end;

architecture behav of tb is
begin
  assert false report "end" severity note;
end behav;
