
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2415.vhd,v 1.2 2001-10-26 16:29:47 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c07s03b02x00p10n01i02415ent IS
END c07s03b02x00p10n01i02415ent;

ARCHITECTURE c07s03b02x00p10n01i02415arch OF c07s03b02x00p10n01i02415ent IS
  type sigrec1 is
    record
      B1 : bit;
      B2 : integer;
      B3 : bit;
    end record;
  
  signal S1 : bit;
  signal S2 : integer;
  signal S3 : bit;
BEGIN
  TESTING: PROCESS
  BEGIN
    (S1, S2, S3) <= sigrec1'('0', 2, '1');
    wait for 1 ns;
    assert NOT(S1='0' and S2=2 and S3='1')
      report "***PASSED TEST: c07s03b02x00p10n01i02415" 
      severity NOTE;
    assert (S1='0' and S2=2 and S3='1')
      report "***FAILED TEST: c07s03b02x00p10n01i02415 - Type of the aggregate must be determinable from the context."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c07s03b02x00p10n01i02415arch;
