
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1423.vhd,v 1.2 2001-10-26 16:29:41 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c08s06b00x00p05n01i01423ent IS
END c08s06b00x00p05n01i01423ent;

ARCHITECTURE c08s06b00x00p05n01i01423arch OF c08s06b00x00p05n01i01423ent IS
  procedure check (signal x   : in  integer;
                   signal kkk : out integer ) is
  begin
    if (x = 0) then
      kkk <= 5;
      wait for 1 ns;
    end if;
  end check;
  signal k  : integer := 0;
  signal kk  : integer := 0;
BEGIN
  TESTING : PROCESS
  BEGIN
    check (k,kk);
    assert NOT(kk = 5)
      report "***PASSED TEST: c08s06b00x00p05n01i01423"
      severity NOTE;
    assert (kk = 5)
      report "***FAILED TEST: c08s06b00x00p05n01i01423 - No actual parmeter is required for a formal parmeter with a default expression."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c08s06b00x00p05n01i01423arch;
