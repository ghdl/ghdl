package pkg is
  constant a : integer := 5; -- Strange but valid character: é
  --  Invalid ascii character 
end pkg;
