entity a is
  constant c : natural := std'u;
end;
