package pkgb is
  shared variable v : natural;
end pkgb;
