library ieee;
use ieee.std_logic_1164.all;

entity t2 is
end t2;

architecture behav of t2 is
  constant my_const : std_ulogic_vector := "01XWL";
  constant my_str : string := "Hello";
begin
end;
