architecturerestrict[=to 0