library ieee;use ieee.std_logic_1164;entity ghdlcrash is
port(i:std'l);end ghdlcrash;architecture s of h is--
function m(a:l)return n is
variable m:t;begin--
end function;--
begin--
end architecture;