configuration"
"
for