entity repro1 is
end;

architecture behav of repro1 is
  constant c : natural := 5 % 4;
begin
end;
