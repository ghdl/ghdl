
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library std;
use std.textio.all;

entity tb is
end tb;

architecture augh of tb is

	constant simu_max_cycles : natural := 1000000;
	constant simu_disp_cycles : std_logic := '0';
	constant simu_err_end_in : std_logic := '0';
	constant reset_cycles : natural := 4;

	component top is
		port (
			clock : in  std_logic;
			reset : in  std_logic;
			start : in  std_logic;
			stdout_rdy : out std_logic;
			stdout_ack : in  std_logic;
			stdin_ack : in  std_logic;
			stdout_data : out std_logic_vector(7 downto 0);
			stdin_data : in  std_logic_vector(7 downto 0);
			stdin_rdy : out std_logic
		);
	end component;

	signal clock : std_logic := '0';
	signal reset : std_logic := '0';
	signal start : std_logic := '0';

	signal clock_next : std_logic := '0';

	-- Access 'clock' model 'clock'

	-- Access 'reset' model 'reset'

	-- Access 'start' model 'start'

	-- Access 'stdin' model 'fifo_in'
	signal stdin_data : std_logic_vector(7 downto 0) := (others => '0');
	signal stdin_rdy : std_logic := '0';
	signal stdin_ack : std_logic := '0';
	signal stdin_vector_idx : natural := 0;
	signal stdin_vector : std_logic_vector(7 downto 0) := (others => '0');
	-- Test vectors
	constant stdin_vectors_nb : natural := 5207;
	type stdin_vec_type is array (0 to stdin_vectors_nb-1) of std_logic_vector(7 downto 0);
	constant stdin_vectors : stdin_vec_type := (
		X"ff", X"d8", X"ff", X"e0", X"00", X"10", X"4a", X"46", X"49", X"46", X"00", X"01", X"01", X"00", X"00",
		X"01", X"00", X"01", X"00", X"00", X"ff", X"db", X"00", X"43", X"00", X"03", X"02", X"02", X"02", X"02",
		X"02", X"03", X"02", X"02", X"02", X"03", X"03", X"03", X"03", X"04", X"06", X"04", X"04", X"04", X"04",
		X"04", X"08", X"06", X"06", X"05", X"06", X"09", X"08", X"0a", X"0a", X"09", X"08", X"09", X"09", X"0a",
		X"0c", X"0f", X"0c", X"0a", X"0b", X"0e", X"0b", X"09", X"09", X"0d", X"11", X"0d", X"0e", X"0f", X"10",
		X"10", X"11", X"10", X"0a", X"0c", X"12", X"13", X"12", X"10", X"13", X"0f", X"10", X"10", X"10", X"ff",
		X"db", X"00", X"43", X"01", X"03", X"03", X"03", X"04", X"03", X"04", X"08", X"04", X"04", X"08", X"10",
		X"0b", X"09", X"0b", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10",
		X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10",
		X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10",
		X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"10", X"ff", X"c0", X"00", X"11", X"08", X"00", X"3b",
		X"00", X"5a", X"03", X"01", X"22", X"00", X"02", X"11", X"01", X"03", X"11", X"01", X"ff", X"c4", X"00",
		X"1f", X"00", X"00", X"01", X"05", X"01", X"01", X"01", X"01", X"01", X"01", X"00", X"00", X"00", X"00",
		X"00", X"00", X"00", X"00", X"01", X"02", X"03", X"04", X"05", X"06", X"07", X"08", X"09", X"0a", X"0b",
		X"ff", X"c4", X"00", X"b5", X"10", X"00", X"02", X"01", X"03", X"03", X"02", X"04", X"03", X"05", X"05",
		X"04", X"04", X"00", X"00", X"01", X"7d", X"01", X"02", X"03", X"00", X"04", X"11", X"05", X"12", X"21",
		X"31", X"41", X"06", X"13", X"51", X"61", X"07", X"22", X"71", X"14", X"32", X"81", X"91", X"a1", X"08",
		X"23", X"42", X"b1", X"c1", X"15", X"52", X"d1", X"f0", X"24", X"33", X"62", X"72", X"82", X"09", X"0a",
		X"16", X"17", X"18", X"19", X"1a", X"25", X"26", X"27", X"28", X"29", X"2a", X"34", X"35", X"36", X"37",
		X"38", X"39", X"3a", X"43", X"44", X"45", X"46", X"47", X"48", X"49", X"4a", X"53", X"54", X"55", X"56",
		X"57", X"58", X"59", X"5a", X"63", X"64", X"65", X"66", X"67", X"68", X"69", X"6a", X"73", X"74", X"75",
		X"76", X"77", X"78", X"79", X"7a", X"83", X"84", X"85", X"86", X"87", X"88", X"89", X"8a", X"92", X"93",
		X"94", X"95", X"96", X"97", X"98", X"99", X"9a", X"a2", X"a3", X"a4", X"a5", X"a6", X"a7", X"a8", X"a9",
		X"aa", X"b2", X"b3", X"b4", X"b5", X"b6", X"b7", X"b8", X"b9", X"ba", X"c2", X"c3", X"c4", X"c5", X"c6",
		X"c7", X"c8", X"c9", X"ca", X"d2", X"d3", X"d4", X"d5", X"d6", X"d7", X"d8", X"d9", X"da", X"e1", X"e2",
		X"e3", X"e4", X"e5", X"e6", X"e7", X"e8", X"e9", X"ea", X"f1", X"f2", X"f3", X"f4", X"f5", X"f6", X"f7",
		X"f8", X"f9", X"fa", X"ff", X"c4", X"00", X"1f", X"01", X"00", X"03", X"01", X"01", X"01", X"01", X"01",
		X"01", X"01", X"01", X"01", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"02", X"03", X"04", X"05",
		X"06", X"07", X"08", X"09", X"0a", X"0b", X"ff", X"c4", X"00", X"b5", X"11", X"00", X"02", X"01", X"02",
		X"04", X"04", X"03", X"04", X"07", X"05", X"04", X"04", X"00", X"01", X"02", X"77", X"00", X"01", X"02",
		X"03", X"11", X"04", X"05", X"21", X"31", X"06", X"12", X"41", X"51", X"07", X"61", X"71", X"13", X"22",
		X"32", X"81", X"08", X"14", X"42", X"91", X"a1", X"b1", X"c1", X"09", X"23", X"33", X"52", X"f0", X"15",
		X"62", X"72", X"d1", X"0a", X"16", X"24", X"34", X"e1", X"25", X"f1", X"17", X"18", X"19", X"1a", X"26",
		X"27", X"28", X"29", X"2a", X"35", X"36", X"37", X"38", X"39", X"3a", X"43", X"44", X"45", X"46", X"47",
		X"48", X"49", X"4a", X"53", X"54", X"55", X"56", X"57", X"58", X"59", X"5a", X"63", X"64", X"65", X"66",
		X"67", X"68", X"69", X"6a", X"73", X"74", X"75", X"76", X"77", X"78", X"79", X"7a", X"82", X"83", X"84",
		X"85", X"86", X"87", X"88", X"89", X"8a", X"92", X"93", X"94", X"95", X"96", X"97", X"98", X"99", X"9a",
		X"a2", X"a3", X"a4", X"a5", X"a6", X"a7", X"a8", X"a9", X"aa", X"b2", X"b3", X"b4", X"b5", X"b6", X"b7",
		X"b8", X"b9", X"ba", X"c2", X"c3", X"c4", X"c5", X"c6", X"c7", X"c8", X"c9", X"ca", X"d2", X"d3", X"d4",
		X"d5", X"d6", X"d7", X"d8", X"d9", X"da", X"e2", X"e3", X"e4", X"e5", X"e6", X"e7", X"e8", X"e9", X"ea",
		X"f2", X"f3", X"f4", X"f5", X"f6", X"f7", X"f8", X"f9", X"fa", X"ff", X"da", X"00", X"0c", X"03", X"01",
		X"00", X"02", X"11", X"03", X"11", X"00", X"3f", X"00", X"f5", X"af", X"00", X"5a", X"ea", X"17", X"b3",
		X"af", X"8a", X"3c", X"4f", X"31", X"f1", X"a4", X"7a", X"9b", X"cf", X"a9", X"e9", X"be", X"22", X"b0",
		X"67", X"16", X"7a", X"6c", X"56", X"f1", X"2a", X"5b", X"da", X"ac", X"0c", X"49", X"2c", X"c7", X"cc",
		X"26", X"40", X"19", X"64", X"2c", X"78", X"e3", X"0b", X"c0", X"e8", X"ba", X"37", X"ed", X"3b", X"a3",
		X"4d", X"e3", X"4d", X"3b", X"5b", X"f1", X"7f", X"85", X"35", X"4d", X"06", X"d2", X"d6", X"e2", X"f6",
		X"3b", X"b8", X"44", X"f0", X"dd", X"58", X"4b", X"72", X"04", X"88", X"33", X"90", X"56", X"28", X"90",
		X"3c", X"98", X"2c", X"55", X"be", X"51", X"ec", X"bf", X"2a", X"78", X"33", X"f6", X"8b", X"f1", X"0f",
		X"c2", X"5f", X"88", X"6d", X"a4", X"45", X"ac", X"ea", X"67", X"c2", X"d1", X"de", X"2c", X"71", X"da",
		X"c3", X"75", X"98", X"23", X"b6", X"91", X"8c", X"8c", X"21", X"8d", X"b7", X"04", X"43", X"bf", X"20",
		X"20", X"00", X"02", X"70", X"3a", X"57", X"b0", X"f8", X"17", X"f6", X"c6", X"f0", X"c0", X"f1", X"61",
		X"f1", X"47", X"88", X"fc", X"31", X"2c", X"1a", X"bf", X"8e", X"ae", X"23", X"b6", X"ba", X"d5", X"12",
		X"ff", X"00", X"cb", X"b6", X"d2", X"74", X"f5", X"8e", X"3b", X"68", X"a4", X"72", X"dc", X"c8", X"04",
		X"b0", X"b3", X"48", X"59", X"40", X"0a", X"c4", X"8e", X"a5", X"1f", X"b7", X"0d", X"8e", X"a5", X"cf",
		X"19", X"29", X"6b", X"36", X"9b", X"be", X"9a", X"35", X"b7", X"9e", X"bd", X"fe", X"f3", X"17", X"24",
		X"d2", X"e8", X"7d", X"0b", X"a9", X"6a", X"16", X"1e", X"35", X"f8", X"18", X"26", X"f1", X"4e", X"81",
		X"a4", X"78", X"96", X"4d", X"46", X"da", X"3b", X"e9", X"2d", X"74", X"eb", X"69", X"ef", X"ed", X"75",
		X"0b", X"79", X"44", X"5b", X"af", X"e3", X"8a", X"75", X"8e", X"48", X"90", X"0d", X"d3", X"18", X"93",
		X"2c", X"81", X"41", X"52", X"e1", X"81", X"3f", X"28", X"f8", X"93", X"f6", X"61", X"f0", X"ab", X"93",
		X"a6", X"e8", X"cf", X"ac", X"4b", X"7f", X"73", X"31", X"6b", X"3b", X"ab", X"0b", X"79", X"2f", X"74",
		X"bb", X"a8", X"e5", X"5d", X"e9", X"11", X"5c", X"97", X"b7", X"75", X"1f", X"2e", X"72", X"c1", X"80",
		X"1d", X"49", X"c0", X"fa", X"ab", X"c5", X"9e", X"0a", X"ba", X"d7", X"be", X"c9", X"1b", X"f8", X"aa",
		X"d6", X"ee", X"41", X"63", X"75", X"35", X"be", X"95", X"67", X"6b", X"1d", X"c5", X"94", X"93", X"88",
		X"d5", X"33", X"05", X"c7", X"dd", X"b7", X"3c", X"43", X"22", X"92", X"e1", X"88", X"32", X"2f", X"28",
		X"5e", X"bc", X"27", X"e1", X"87", X"c5", X"4f", X"8c", X"b0", X"7c", X"47", X"82", X"d3", X"c4", X"63",
		X"56", X"9f", X"45", X"b4", X"69", X"2d", X"66", X"d2", X"ac", X"6d", X"12", X"5b", X"95", X"73", X"84",
		X"86", X"6d", X"eb", X"f2", X"ac", X"46", X"56", X"60", X"1d", X"9f", X"0e", X"55", X"8f", X"40", X"71",
		X"ea", X"ca", X"18", X"5a", X"8b", X"92", X"b2", X"4d", X"6c", X"b4", X"f4", X"d2", X"fd", X"1d", X"ff",
		X"00", X"22", X"bc", X"d9", X"f3", X"4f", X"c2", X"cd", X"43", X"c7", X"1f", X"03", X"be", X"25", X"e9",
		X"5e", X"2b", X"83", X"45", X"7d", X"28", X"43", X"a8", X"bf", X"87", X"ef", X"6e", X"ae", X"ad", X"9f",
		X"ec", X"f1", X"c9", X"24", X"8a", X"b2", X"c5", X"b9", X"86", X"03", X"aa", X"ec", X"6f", X"50", X"3b",
		X"57", X"d6", X"1f", X"b5", X"64", X"2b", X"60", X"9a", X"45", X"97", X"88", X"fc", X"09", X"a0", X"9b",
		X"5d", X"50", X"c5", X"a8", X"b6", X"a5", X"16", X"9e", X"0c", X"df", X"68", X"52", X"43", X"42", X"d2",
		X"e0", X"61", X"f2", X"01", X"20", X"9e", X"47", X"6e", X"e3", X"63", X"e1", X"6f", X"c3", X"2f", X"09",
		X"7c", X"45", X"b6", X"f1", X"2f", X"8a", X"7c", X"75", X"3e", X"bf", X"6e", X"d6", X"7e", X"36", X"d7",
		X"e6", X"b8", X"85", X"54", X"ba", X"31", X"69", X"96", X"23", X"94", X"19", X"8d", X"dc", X"28", X"64",
		X"25", X"79", X"04", X"b1", X"07", X"1c", X"8e", X"b7", X"c3", X"fe", X"28", X"5d", X"41", X"6d", X"3e",
		X"0a", X"7c", X"4a", X"b5", X"d4", X"b5", X"d3", X"a9", X"d9", X"df", X"ed", X"d4", X"2e", X"ed", X"a1",
		X"31", X"6a", X"91", X"c5", X"b5", X"44", X"de", X"64", X"60", X"20", X"66", X"59", X"10", X"02", X"83",
		X"76", X"76", X"93", X"8e", X"b5", X"e7", X"52", X"c0", X"ca", X"ae", X"0e", X"58", X"6a", X"53", X"b7",
		X"3a", X"de", X"d7", X"b5", X"fa", X"7c", X"cc", X"b5", X"94", X"4f", X"84", X"3c", X"49", X"06", X"b3",
		X"ac", X"47", X"7d", X"ab", X"5c", X"da", X"ac", X"96", X"92", X"30", X"36", X"a8", X"17", X"e4", X"b7",
		X"80", X"1c", X"02", X"3d", X"73", X"ec", X"3b", X"f1", X"c5", X"69", X"7c", X"21", X"f8", X"07", X"e2",
		X"af", X"8e", X"1a", X"f3", X"be", X"9d", X"ac", X"db", X"da", X"c3", X"a4", X"5f", X"5a", X"a6", X"a1",
		X"6e", X"08", X"37", X"11", X"d9", X"49", X"9f", X"df", X"44", X"87", X"87", X"3b", X"94", X"a6", X"de",
		X"c4", X"e7", X"9c", X"60", X"fd", X"11", X"f1", X"13", X"e0", X"9f", X"82", X"3c", X"2f", X"e1", X"f7",
		X"f0", X"57", X"87", X"6d", X"ae", X"13", X"59", X"f0", X"ed", X"bc", X"7a", X"c5", X"ad", X"c5", X"c9",
		X"95", X"ee", X"1b", X"4f", X"09", X"fb", X"d5", X"b8", X"91", X"9b", X"cb", X"7e", X"59", X"86", X"11",
		X"72", X"18", X"02", X"00", X"c1", X"af", X"09", X"f8", X"7d", X"e1", X"6f", X"88", X"56", X"9e", X"3b",
		X"8f", X"e2", X"0f", X"c2", X"2d", X"40", X"4b", X"3c", X"12", X"ad", X"ac", X"d0", X"29", X"3e", X"4b",
		X"dc", X"05", X"12", X"24", X"05", X"41", X"07", X"6b", X"0e", X"41", X"cf", X"5e", X"87", X"9c", X"0f",
		X"03", X"0f", X"95", X"d5", X"c1", X"62", X"a1", X"4e", X"b2", X"52", X"4d", X"74", X"76", X"fc", X"ec",
		X"f4", X"ea", X"ec", X"34", X"ef", X"2d", X"74", X"b1", X"ce", X"fc", X"6d", X"f8", X"0b", X"f1", X"13",
		X"e1", X"7f", X"89", X"b5", X"4b", X"7b", X"ab", X"35", X"b9", X"d2", X"22", X"bc", X"5b", X"7d", X"3e",
		X"ea", X"58", X"d6", X"29", X"6f", X"22", X"c2", X"95", X"6d", X"99", X"e0", X"e0", X"95", X"3d", X"06",
		X"53", X"23", X"ae", X"2b", X"99", X"f1", X"77", X"81", X"67", X"9b", X"5b", X"82", X"e6", X"c3", X"4d",
		X"91", X"55", X"ec", X"95", X"b7", X"05", X"c0", X"46", X"f9", X"ba", X"fe", X"95", X"ec", X"3f", X"17",
		X"3e", X"3e", X"f8", X"eb", X"e2", X"b7", X"8a", X"75", X"6f", X"02", X"f8", X"db", X"51", X"b7", X"d1",
		X"6f", X"6d", X"8a", X"db", X"c3", X"6b", X"0c", X"2a", X"b1", X"f9", X"e8", X"a0", X"ed", X"67", X"70",
		X"64", X"ce", X"7d", X"ff", X"00", X"a8", X"a6", X"7c", X"2e", X"b6", X"f1", X"ce", X"b1", X"e1", X"7b",
		X"cb", X"1f", X"16", X"e8", X"b3", X"33", X"08", X"64", X"fb", X"2d", X"d2", X"5b", X"b3", X"29", X"74",
		X"18", X"20", X"b0", X"18", X"ef", X"eb", X"5e", X"66", X"73", X"56", X"50", X"c5", X"3f", X"ab", X"a7",
		X"ee", X"e8", X"d3", X"f3", X"fc", X"d7", X"99", X"a2", X"69", X"e8", X"d9", X"f3", X"76", X"9b", X"6d",
		X"a8", X"68", X"b7", X"d1", X"dd", X"6a", X"9a", X"44", X"b3", X"24", X"33", X"6e", X"90", X"94", X"3b",
		X"5b", X"19", X"f5", X"ea", X"2b", X"aa", X"7f", X"11", X"f8", X"76", X"57", X"69", X"17", X"45", X"da",
		X"1c", X"96", X"03", X"6a", X"f0", X"0f", X"e3", X"51", X"6a", X"ba", X"37", X"8c", X"5b", X"75", X"f5",
		X"d5", X"b5", X"cb", X"da", X"29", X"2c", X"e2", X"3c", X"10", X"07", X"51", X"90", X"39", X"ee", X"3f",
		X"ad", X"72", X"0f", X"1d", X"e1", X"76", X"29", X"6d", X"31", X"52", X"4e", X"38", X"23", X"8a", X"ba",
		X"78", X"87", X"6b", X"e8", X"5f", X"3b", X"a7", X"a2", X"47", X"af", X"fc", X"24", X"f8", X"75", X"17",
		X"8e", X"6e", X"af", X"6f", X"f5", X"dd", X"5b", X"4b", X"83", X"4f", X"b3", X"b8", X"d2", X"ac", X"5e",
		X"39", X"e4", X"58", X"6f", X"24", X"8a", X"e2", X"ee", X"18", X"44", X"d6", X"ca", X"e3", X"1b", X"11",
		X"58", X"a3", X"15", X"63", X"b0", X"b4", X"7d", X"b1", X"9f", X"4c", X"f8", X"a1", X"fb", X"3f", X"4d",
		X"f0", X"ef", X"c1", X"56", X"97", X"fa", X"c6", X"89", X"f6", X"bd", X"13", X"53", X"b3", X"3f", X"d8",
		X"ba", X"ea", X"98", X"18", X"3a", X"cd", X"03", X"4d", X"f6", X"79", X"c0", X"61", X"22", X"31", X"c6",
		X"e5", X"23", X"31", X"b9", X"73", X"80", X"4b", X"28", X"ae", X"2b", X"e1", X"bf", X"c4", X"8d", X"5b",
		X"e0", X"67", X"ed", X"10", X"fe", X"13", X"f0", X"d6", X"a6", X"97", X"5e", X"16", X"83", X"56", X"1a",
		X"72", X"3f", X"88", X"a5", X"fb", X"27", X"d9", X"2c", X"ae", X"1e", X"30", X"f2", X"79", X"b2", X"30",
		X"5b", X"60", X"aa", X"cc", X"cc", X"dc", X"23", X"a2", X"7c", X"c3", X"a1", X"1f", X"50", X"7c", X"46",
		X"f1", X"ee", X"81", X"e3", X"4d", X"63", X"e2", X"2e", X"91", X"e1", X"bd", X"6f", X"43", X"d4", X"fc",
		X"05", X"a0", X"f8", X"6a", X"35", X"36", X"f1", X"5f", X"db", X"cd", X"61", X"79", X"af", X"dd", X"c3",
		X"21", X"86", X"4b", X"49", X"1c", X"c8", X"b1", X"a5", X"bc", X"2c", X"f3", X"4a", X"b1", X"15", X"5f",
		X"b5", X"30", X"0f", X"b5", X"d0", X"4d", X"5f", X"4b", X"83", X"8e", X"1e", X"78", X"58", X"ca", X"1a",
		X"bb", X"3e", X"8b", X"aa", X"6f", X"ce", X"eb", X"5f", X"91", X"ce", X"e1", X"6b", X"a7", X"b8", X"bf",
		X"09", X"35", X"5f", X"88", X"5e", X"29", X"b0", X"f0", X"96", X"a1", X"f1", X"93", X"5a", X"7d", X"57",
		X"4c", X"f1", X"4e", X"99", X"35", X"c8", X"b1", X"93", X"58", X"5b", X"78", X"e3", X"d3", X"e1", X"b6",
		X"1e", X"5d", X"e1", X"59", X"08", X"59", X"1c", X"80", X"b1", X"ba", X"e1", X"54", X"2c", X"8d", X"b9",
		X"c3", X"90", X"6b", X"85", X"f1", X"3f", X"83", X"fc", X"2d", X"e1", X"4f", X"07", X"fc", X"5d", X"d5",
		X"fe", X"19", X"fc", X"6e", X"bb", X"d4", X"7c", X"29", X"a4", X"5b", X"a3", X"c9", X"a5", X"41", X"a5",
		X"bd", X"f4", X"f1", X"86", X"8d", X"02", X"b4", X"17", X"30", X"4c", X"82", X"35", X"f3", X"83", X"c4",
		X"66", X"75", X"61", X"09", X"8c", X"97", X"69", X"4f", X"cd", X"5e", X"25", X"e0", X"ff", X"00", X"da",
		X"03", X"e2", X"87", X"84", X"ed", X"cc", X"9a", X"6e", X"af", X"0c", X"49", X"e1", X"bd", X"1e", X"ff",
		X"00", X"c3", X"16", X"8b", X"3d", X"a2", X"c8", X"23", X"b5", X"bc", X"1b", X"c6", X"c0", X"c5", X"70",
		X"c2", X"65", X"50", X"c5", X"9b", X"05", X"42", X"8c", X"65", X"4a", X"bf", X"d8", X"bf", X"00", X"61",
		X"f8", X"6a", X"9e", X"11", X"f0", X"d6", X"9d", X"e2", X"4d", X"1f", X"c3", X"1a", X"6e", X"b3", X"a6",
		X"da", X"47", X"a4", X"a0", X"b3", X"d7", X"ad", X"22", X"96", X"7b", X"50", X"88", X"d0", X"a4", X"72",
		X"cf", X"2c", X"72", X"2c", X"b2", X"0f", X"20", X"14", X"24", X"6f", X"95", X"37", X"2b", X"48", X"85",
		X"56", X"2d", X"b0", X"53", X"86", X"63", X"15", X"da", X"1b", X"b6", X"9d", X"f5", X"5b", X"5d", X"5b",
		X"c9", X"ef", X"aa", X"dc", X"77", X"ba", X"b9", X"f3", X"af", X"ec", X"cd", X"f1", X"73", X"54", X"d3",
		X"3c", X"4b", X"e2", X"af", X"0c", X"cd", X"e1", X"0d", X"0a", X"fe", X"43", X"e1", X"8d", X"4f", X"53",
		X"b6", X"d6", X"67", X"d2", X"fc", X"eb", X"bb", X"1b", X"b7", X"b2", X"31", X"ed", X"92", X"6c", X"11",
		X"24", X"77", X"12", X"98", X"d5", X"84", X"d8", X"05", X"c0", X"c3", X"1c", X"98", X"64", X"f5", X"ef",
		X"8b", X"1f", X"17", X"bc", X"2d", X"a5", X"78", X"a7", X"c0", X"9e", X"2c", X"bc", X"d2", X"75", X"3f",
		X"0d", X"78", X"4e", X"e8", X"8d", X"5b", X"49", X"f1", X"6e", X"9f", X"6c", X"d2", X"4b", X"67", X"6c",
		X"61", X"49", X"a1", X"d3", X"84", X"20", X"b4", X"4e", X"a1", X"27", X"41", X"36", X"e4", X"95", X"c8",
		X"56", X"55", X"89", X"3e", X"fa", X"75", X"df", X"13", X"7e", X"1b", X"68", X"5f", X"0b", X"7e", X"1d",
		X"cd", X"ab", X"7c", X"1a", X"9f", X"48", X"16", X"f0", X"de", X"dd", X"e8", X"fe", X"27", X"68", X"a4",
		X"82", X"e2", X"7d", X"52", X"01", X"20", X"2e", X"cf", X"1c", X"5f", X"bb", X"17", X"51", X"f9", X"9b",
		X"37", X"48", X"81", X"a3", X"42", X"a2", X"3f", X"2f", X"e4", X"65", X"e1", X"ac", X"be", X"20", X"78",
		X"93", X"4a", X"fd", X"9d", X"fc", X"21", X"e1", X"7f", X"08", X"78", X"72", X"e2", X"0d", X"4e", X"e6",
		X"4b", X"9b", X"09", X"75", X"b9", X"46", X"fb", X"3b", X"6b", X"bb", X"59", X"96", X"d7", X"ce", X"5d",
		X"e1", X"97", X"73", X"47", X"22", X"c2", X"61", X"0a", X"a5", X"9f", X"2d", X"b7", X"6a", X"c8", X"e1",
		X"61", X"e7", X"57", X"0d", X"28", X"51", X"a5", X"53", X"9b", X"dd", X"be", X"9e", X"4d", X"2d", X"15",
		X"fe", X"57", X"d0", X"13", X"e5", X"f7", X"64", X"b5", X"47", X"b4", X"bf", X"8a", X"be", X"1c", X"7c",
		X"61", X"f0", X"a6", X"a6", X"da", X"6e", X"a3", X"e1", X"3f", X"17", X"e2", X"c2", X"56", X"d2", X"ed",
		X"6d", X"23", X"b8", X"d2", X"b5", X"18", X"6f", X"17", X"ce", X"8e", X"7f", X"31", X"26", X"67", X"68",
		X"c4", X"cc", X"47", X"96", X"ee", X"9b", X"4a", X"c8", X"bb", X"81", X"18", X"91", X"be", X"78", X"f8",
		X"51", X"1e", X"b1", X"f0", X"33", X"c4", X"f1", X"f8", X"a2", X"3f", X"0e", X"1f", X"15", X"e8", X"9e",
		X"3c", X"10", X"be", X"92", X"d1", X"c5", X"2d", X"b4", X"6b", X"22", X"39", X"60", X"e8", X"85", X"49",
		X"f9", X"06", X"ec", X"b9", X"00", X"61", X"41", X"ca", X"f7", X"e0", X"bc", X"59", X"e3", X"7d", X"4f",
		X"c4", X"3e", X"1f", X"f0", X"50", X"f8", X"68", X"b6", X"b6", X"7a", X"a4", X"fa", X"79", X"b7", X"d4",
		X"35", X"4b", X"6d", X"3e", X"0b", X"09", X"2c", X"2e", X"2d", X"94", X"5b", X"0b", X"51", X"2c", X"67",
		X"76", X"c5", X"8d", X"0c", X"68", X"32", X"59", X"91", X"57", X"92", X"0e", X"17", X"d9", X"fe", X"16",
		X"fc", X"5c", X"d4", X"fe", X"25", X"69", X"3e", X"09", X"f0", X"3f", X"c6", X"af", X"14", X"58", X"69",
		X"16", X"ba", X"ad", X"dd", X"ed", X"c4", X"17", X"2d", X"1a", X"c1", X"3e", X"bb", X"24", X"8d", X"24",
		X"96", X"ca", X"e5", X"00", X"55", X"59", X"da", X"48", X"f0", X"aa", X"23", X"59", X"54", X"c2", X"18",
		X"16", X"68", X"98", X"63", X"88", X"cc", X"69", X"54", X"94", X"53", X"4f", X"9a", X"fa", X"3f", X"37",
		X"6d", X"35", X"ec", X"9b", X"ba", X"7b", X"7c", X"8b", X"94", X"5a", X"d5", X"1e", X"5b", X"f1", X"bf",
		X"c0", X"e3", X"c6", X"3f", X"1d", X"63", X"f1", X"57", X"8c", X"fc", X"3d", X"ab", X"6a", X"1e", X"10",
		X"b5", X"45", X"b8", X"9b", X"4a", X"d3", X"9a", X"2b", X"7b", X"d8", X"92", X"4d", X"a2", X"49", X"96",
		X"68", X"f1", X"e6", X"95", X"25", X"18", X"82", X"41", X"23", X"1e", X"a0", X"1f", X"a3", X"93", X"5b",
		X"d0", X"3f", X"67", X"3d", X"36", X"d2", X"18", X"35", X"1d", X"74", X"f8", X"56", X"dd", X"63", X"b7",
		X"bb", X"63", X"7a", X"93", X"35", X"bd", X"c3", X"8d", X"f0", X"0c", X"9c", X"b6", X"46", X"c6", X"dc",
		X"31", X"b4", X"ef", X"03", X"3c", X"f1", X"f2", X"8f", X"c5", X"7d", X"7f", X"c6", X"bf", X"0e", X"3c",
		X"63", X"af", X"78", X"20", X"6b", X"8e", X"9a", X"cc", X"16", X"e8", X"2f", X"05", X"cc", X"6a", X"ef",
		X"77", X"1c", X"cb", X"e6", X"b8", X"ca", X"91", X"1a", X"60", X"30", X"04", X"2e", X"39", X"c0", X"18",
		X"0a", X"b4", X"db", X"9d", X"1f", X"c5", X"91", X"fc", X"1a", X"b7", X"d7", X"ae", X"7e", X"d6", X"ba",
		X"1f", X"89", X"6d", X"a3", X"32", X"dd", X"5c", X"93", X"3c", X"6c", X"d1", X"b9", X"75", X"d8", X"d9",
		X"26", X"26", X"0c", X"a4", X"15", X"eb", X"80", X"78", X"ca", X"a8", X"3c", X"f5", X"f3", X"08", X"c2",
		X"53", X"53", X"83", X"72", X"57", X"bf", X"5b", X"2e", X"97", X"6b", X"a6", X"da", X"8d", X"2d", X"39",
		X"91", X"8b", X"fb", X"45", X"eb", X"7f", X"08", X"64", X"d6", X"66", X"f1", X"0f", X"c1", X"8d", X"46",
		X"45", X"8f", X"57", X"bb", X"37", X"32", X"5a", X"01", X"32", X"47", X"6a", X"c7", X"e6", X"90", X"04",
		X"93", X"3b", X"54", X"b9", X"61", X"b0", X"70", X"0e", X"ec", X"71", X"8a", X"e2", X"ad", X"f5", X"4d",
		X"2d", X"e0", X"8d", X"e7", X"4b", X"33", X"2b", X"20", X"2e", X"41", X"1f", X"7b", X"1c", X"fe", X"b5",
		X"cd", X"d8", X"e8", X"76", X"fa", X"cc", X"1a", X"84", X"cf", X"2b", X"46", X"22", X"96", X"35", X"0e",
		X"4f", X"0a", X"a5", X"b0", X"c4", X"8f", X"a6", X"33", X"5d", X"3a", X"f8", X"23", X"c1", X"b1", X"01",
		X"19", X"f1", X"cd", X"be", X"50", X"6d", X"e0", X"8c", X"71", X"5f", X"35", X"88", X"9d", X"1c", X"44",
		X"dc", X"9a", X"e5", X"f2", X"5f", X"d3", X"1c", X"6a", X"24", X"bd", X"e4", X"68", X"78", X"8b", X"44",
		X"f0", X"ec", X"da", X"fe", X"bd", X"af", X"db", X"c7", X"7d", X"76", X"fa", X"14", X"33", X"d9", X"6a",
		X"36", X"80", X"2c", X"72", X"c1", X"3b", X"20", X"84", X"5d", X"c6", X"1c", X"62", X"48", X"c5", X"c3",
		X"10", X"f1", X"fc", X"ad", X"1c", X"8f", X"b8", X"36", X"d9", X"03", X"2f", X"a7", X"ff", X"00", X"c3",
		X"33", X"fc", X"67", X"f0", X"b7", X"84", X"2d", X"b4", X"81", X"af", X"46", X"3c", X"0b", X"af", X"db",
		X"db", X"6b", X"17", X"d7", X"30", X"44", X"b7", X"36", X"31", X"7d", X"a6", X"28", X"51", X"ae", X"15",
		X"23", X"6f", X"32", X"e3", X"74", X"2d", X"1c", X"70", X"be", X"e8", X"c7", X"ef", X"48", X"dc", X"8c",
		X"ec", X"4f", X"55", X"f0", X"9b", X"c0", X"5e", X"24", X"f8", X"ef", X"e3", X"73", X"e2", X"3f", X"8a",
		X"de", X"0f", X"d2", X"bc", X"67", X"e1", X"d1", X"a7", X"5a", X"e9", X"57", X"da", X"9f", X"9f", X"71",
		X"63", X"a9", X"d8", X"8b", X"76", X"91", X"62", X"b9", X"83", X"0c", X"66", X"95", X"d1", X"da", X"48",
		X"4b", X"30", X"c9", X"8a", X"dd", X"17", X"92", X"be", X"5b", X"7d", X"57", X"a9", X"dd", X"7c", X"3d",
		X"d0", X"74", X"25", X"f1", X"26", X"9f", X"71", X"ac", X"7d", X"8f", X"e1", X"d6", X"b5", X"a9", X"59",
		X"bd", X"b6", X"96", X"a2", X"ce", X"0b", X"78", X"84", X"9b", X"2f", X"8d", X"ea", X"a1", X"2b", X"39",
		X"42", X"af", X"bb", X"04", X"0c", X"dc", X"b1", X"95", X"76", X"3b", X"13", X"f4", X"58", X"5c", X"05",
		X"e3", X"2a", X"94", X"fd", X"e8", X"b7", X"a5", X"9d", X"b4", X"4f", X"55", X"d9", X"ad", X"f6", X"ec",
		X"65", X"0f", X"79", X"dd", X"bb", X"1f", X"9d", X"ba", X"97", X"86", X"f4", X"af", X"0f", X"fc", X"6f",
		X"d6", X"fc", X"31", X"6d", X"e2", X"4b", X"58", X"b4", X"6d", X"33", X"56", X"2e", X"d7", X"9a", X"b5",
		X"a1", X"78", X"a6", X"8e", X"39", X"be", X"d1", X"e6", X"cb", X"6e", X"84", X"99", X"23", X"df", X"13",
		X"6e", X"0a", X"c3", X"f7", X"7b", X"b3", X"91", X"95", X"3c", X"ff", X"00", X"85", X"bc", X"59", X"e1",
		X"2f", X"05", X"78", X"f6", X"df", X"c5", X"2e", X"fa", X"75", X"c5", X"ad", X"b6", X"a3", X"1e", X"a7",
		X"78", X"34", X"dd", X"ab", X"05", X"b4", X"b0", X"dc", X"bb", X"c5", X"1d", X"bc", X"32", X"a3", X"06",
		X"0a", X"c6", X"39", X"55", X"24", X"12", X"21", X"87", X"70", X"71", X"94", X"6c", X"6c", X"7c", X"72",
		X"f8", X"bb", X"73", X"e3", X"2f", X"8a", X"1a", X"cc", X"b6", X"b7", X"16", X"17", X"f6", X"10", X"ea",
		X"da", X"8c", X"b6", X"8d", X"6e", X"64", X"b8", X"b7", X"9d", X"52", X"69", X"13", X"7a", X"97", X"66",
		X"61", X"14", X"d1", X"6e", X"63", X"fc", X"3b", X"5d", X"49", X"1d", X"5a", X"be", X"bf", X"f8", X"11",
		X"63", X"f0", X"5b", X"e2", X"af", X"82", X"fc", X"03", X"a7", X"5e", X"5b", X"6a", X"3a", X"b7", X"88",
		X"fc", X"2a", X"7e", X"cb", X"6b", X"ac", X"6a", X"4a", X"b6", X"ba", X"b5", X"94", X"2b", X"14", X"a0",
		X"b4", X"33", X"08", X"1a", X"29", X"92", X"22", X"1b", X"ca", X"47", X"32", X"15", X"f2", X"b2", X"4b",
		X"bc", X"6a", X"42", X"c0", X"61", X"af", X"5e", X"71", X"a3", X"2d", X"22", X"ee", X"be", X"fb", X"3d",
		X"2f", X"7d", X"3f", X"22", X"69", X"df", X"e1", X"38", X"3f", X"89", X"df", X"b5", X"e7", X"88", X"ad",
		X"7c", X"14", X"9f", X"0f", X"bc", X"15", X"e0", X"af", X"b0", X"78", X"a3", X"5d", X"bf", X"9a", X"f7",
		X"51", X"83", X"54", X"b3", X"33", X"2c", X"fa", X"75", X"d8", X"dd", X"6d", X"76", X"ad", X"03", X"a4",
		X"91", X"5c", X"23", X"14", X"81", X"d6", X"42", X"57", X"71", X"26", X"30", X"ca", X"76", X"47", X"b3",
		X"f0", X"83", X"f6", X"be", X"d1", X"87", X"81", X"63", X"b4", X"f1", X"76", X"ab", X"a7", X"f8", X"7e",
		X"eb", X"46", X"36", X"16", X"b3", X"58", X"59", X"e9", X"41", X"ad", X"f5", X"25", X"78", X"a5", X"8e",
		X"e2", X"f3", X"50", X"88", X"21", X"cc", X"b1", X"4c", X"62", X"90", X"c7", X"a7", X"b4", X"37", X"13",
		X"ca", X"e4", X"ba", X"6c", X"3b", X"e0", X"d1", X"f8", X"45", X"1f", X"c6", X"fb", X"f7", X"f8", X"eb",
		X"f0", X"da", X"f7", X"e1", X"f7", X"85", X"35", X"9f", X"12", X"dc", X"6a", X"0f", X"34", X"96", X"76",
		X"2c", X"5b", X"4d", X"92", X"7b", X"bd", X"38", X"25", X"89", X"33", X"19", X"55", X"e4", X"b6", X"95",
		X"20", X"28", X"9f", X"30", X"65", X"f2", X"e5", X"32", X"fe", X"f0", X"92", X"be", X"35", X"e1", X"bf",
		X"d9", X"e7", X"c5", X"b7", X"82", X"6f", X"05", X"e8", X"b0", X"69", X"7a", X"d6", X"a5", X"76", X"91",
		X"49", X"7f", X"6b", X"7f", X"66", X"22", X"6b", X"4b", X"3d", X"cc", X"b2", X"5e", X"88", X"e4", X"1e",
		X"64", X"8b", X"1c", X"8a", X"b1", X"ae", X"c0", X"ad", X"be", X"64", X"77", X"58", X"95", X"b1", X"5d",
		X"15", X"e1", X"8b", X"a7", X"28", X"fd", X"56", X"f2", X"5b", X"5b", X"6b", X"6b", X"fd", X"6d", X"f9",
		X"1a", X"37", X"ad", X"cb", X"be", X"3f", X"93", X"c2", X"5e", X"20", X"9f", X"5c", X"f0", X"2d", X"b6",
		X"b1", X"75", X"ae", X"69", X"b7", X"9f", X"65", X"6b", X"8f", X"14", X"dd", X"db", X"c9", X"0d", X"d2",
		X"de", X"86", X"50", X"b0", X"a5", X"b9", X"28", X"63", X"91", X"6d", X"62", X"86", X"09", X"8b", X"87",
		X"91", X"76", X"cf", X"08", X"27", X"31", X"ac", X"1e", X"7b", X"a1", X"f8", X"ff", X"00", X"4f", X"d0",
		X"be", X"25", X"5a", X"5d", X"78", X"f3", X"50", X"bb", X"f1", X"46", X"a4", X"b3", X"43", X"69", X"2c",
		X"aa", X"d0", X"25", X"8a", X"69", X"ec", X"88", X"b2", X"43", X"24", X"31", X"29", X"8c", X"6c", X"8d",
		X"42", X"18", X"d0", X"2b", X"2b", X"ab", X"2e", X"55", X"94", X"14", X"e8", X"be", X"12", X"e9", X"16",
		X"13", X"f8", X"8b", X"c3", X"ba", X"a6", X"bd", X"7d", X"77", X"f1", X"17", X"5b", X"d6", X"24", X"6d",
		X"17", X"4a", X"d1", X"2c", X"ee", X"25", X"b4", X"b7", X"96", X"f2", X"65", X"8e", X"d2", X"07", X"b8",
		X"d5", X"2e", X"15", X"45", X"ac", X"42", X"08", X"60", X"2b", X"b0", X"4b", X"23", X"83", X"82", X"10",
		X"39", X"61", X"eb", X"7f", X"0f", X"bf", X"66", X"0f", X"01", X"6b", X"da", X"46", X"9f", X"e3", X"0d",
		X"67", X"c7", X"11", X"f8", X"76", X"da", X"6b", X"fb", X"ab", X"7d", X"62", X"de", X"3d", X"7a", X"d9",
		X"ac", X"6d", X"5a", X"7b", X"b9", X"a0", X"b7", X"f2", X"de", X"45", X"4b", X"88", X"97", X"cf", X"6b",
		X"72", X"ab", X"31", X"de", X"eb", X"21", X"47", X"d9", X"2a", X"18", X"5f", X"9a", X"58", X"6a", X"d9",
		X"8e", X"21", X"d4", X"82", X"49", X"47", X"a3", X"76", X"dd", X"f5", X"7a", X"e9", X"f7", X"bb", X"5c",
		X"6d", X"cd", X"49", X"34", X"70", X"9f", X"b4", X"4c", X"d6", X"df", X"1a", X"34", X"4b", X"7f", X"1d",
		X"f8", X"1e", X"74", X"d5", X"2d", X"34", X"3d", X"3a", X"db", X"51", X"bb", X"8a", X"56", X"8a", X"19",
		X"ed", X"1e", X"67", X"9a", X"27", X"b5", X"44", X"00", X"4f", X"2a", X"2c", X"50", X"a4", X"8e", X"8f",
		X"26", X"e8", X"fc", X"e8", X"88", X"2f", X"92", X"aa", X"9f", X"06", X"ff", X"00", X"69", X"ef", X"86",
		X"f3", X"e9", X"93", X"fc", X"21", X"f8", X"89", X"e1", X"8b", X"58", X"bc", X"3f", X"ac", X"a2", X"5b",
		X"4c", X"ed", X"71", X"04", X"56", X"b0", X"ca", X"54", X"01", X"28", X"8a", X"0b", X"78", X"8c", X"65",
		X"9d", X"e4", X"62", X"e6", X"46", X"23", X"e5", X"0b", X"b7", X"15", X"85", X"f0", X"57", X"c0", X"7a",
		X"cd", X"ff", X"00", X"c4", X"ab", X"9d", X"4d", X"f5", X"4b", X"5b", X"bd", X"17", X"4e", X"bc", X"d4",
		X"34", X"d5", X"8f", X"56", X"bd", X"7b", X"08", X"b5", X"3b", X"74", X"9c", X"c2", X"54", X"4f", X"83",
		X"24", X"8c", X"40", X"24", X"ab", X"23", X"2c", X"60", X"b0", X"28", X"77", X"15", X"af", X"a0", X"fe",
		X"2a", X"7c", X"19", X"f0", X"36", X"a1", X"e2", X"4f", X"16", X"78", X"97", X"c2", X"16", X"da", X"65",
		X"96", X"8f", X"a5", X"68", X"10", X"6a", X"57", X"1a", X"b4", X"d6", X"90", X"b6", X"9f", X"72", X"26",
		X"33", X"ab", X"b5", X"ac", X"fb", X"85", X"bf", X"96", X"be", X"53", X"2c", X"9f", X"bd", X"01", X"1d",
		X"19", X"49", X"db", X"90", X"6a", X"8f", X"b6", X"c5", X"4d", X"d4", X"83", X"49", X"fc", X"2d", X"3d",
		X"53", X"b7", X"45", X"75", X"b7", X"4d", X"cb", X"a7", X"34", X"9d", X"e4", X"ae", X"7c", X"69", X"a2",
		X"d9", X"68", X"3e", X"1f", X"f1", X"c6", X"a3", X"e1", X"9d", X"4b", X"4e", X"b9", X"bc", X"f0", X"a4",
		X"b7", X"93", X"c0", X"93", X"99", X"95", X"84", X"a0", X"33", X"18", X"d0", X"48", X"bc", X"36", X"55",
		X"7d", X"89", X"eb", X"c5", X"74", X"d2", X"f8", X"ab", X"c1", X"91", X"4a", X"f1", X"da", X"7c", X"39",
		X"f0", X"42", X"c0", X"8c", X"56", X"25", X"97", X"51", X"88", X"38", X"40", X"78", X"0c", X"33", X"d7",
		X"18", X"cd", X"72", X"77", X"53", X"68", X"76", X"da", X"65", X"ad", X"87", X"87", X"b5", X"18", X"6f",
		X"d2", X"3d", X"6a", X"62", X"f7", X"a2", X"dd", X"62", X"46", X"90", X"a3", X"32", X"c4", X"02", X"49",
		X"22", X"32", X"8c", X"2a", X"ef", X"56", X"20", X"ef", X"3f", X"dd", X"39", X"e6", X"57", X"e0", X"ac",
		X"5a", X"8a", X"8d", X"41", X"24", X"d5", X"51", X"6e", X"87", X"9c", X"15", X"6c", X"72", X"00", X"6e",
		X"70", X"0e", X"79", X"1c", X"d7", X"cb", X"d5", X"a3", X"05", X"5e", X"71", X"c4", X"3e", X"46", X"9f",
		X"47", X"75", X"bf", X"93", X"35", X"e5", X"e4", X"76", X"86", X"d6", X"4f", X"6b", X"ee", X"77", X"5a",
		X"7f", X"ed", X"43", X"e2", X"cf", X"0e", X"fd", X"a2", X"fb", X"c2", X"7a", X"80", X"d3", X"75", X"3b",
		X"39", X"a3", X"b3", X"5b", X"78", X"96", X"48", X"a1", X"d4", X"34", X"ff", X"00", X"3a", X"39", X"36",
		X"f9", X"8a", X"de", X"6e", X"4c", X"b0", X"a7", X"98", X"85", X"d7", X"7a", X"48", X"fb", X"b7", X"7c",
		X"cb", X"5f", X"5b", X"78", X"eb", X"e2", X"b6", X"bb", X"fb", X"41", X"fc", X"39", X"f1", X"f7", X"86",
		X"24", X"36", X"3e", X"1e", X"d3", X"a7", X"d2", X"b4", X"f5", X"86", X"3b", X"6d", X"5c", X"bd", X"e2",
		X"34", X"86", X"32", X"c8", X"62", X"24", X"33", X"c4", X"b3", X"47", X"2a", X"17", X"09", X"1a", X"6c",
		X"94", X"a9", X"46", X"12", X"b9", X"87", X"f3", X"57", X"c5", X"96", X"d0", X"e9", X"1e", X"28", X"d5",
		X"ec", X"f4", X"e0", X"f1", X"45", X"69", X"ab", X"5c", X"c1", X"0f", X"ce", X"cc", X"ca", X"91", X"ca",
		X"e1", X"06", X"e2", X"49", X"38", X"00", X"72", X"4e", X"78", X"af", X"47", X"f1", X"57", X"8e", X"3c",
		X"4b", X"a3", X"7c", X"28", X"f8", X"69", X"e2", X"cd", X"3e", X"f6", X"14", X"d5", X"a7", X"5d", X"47",
		X"7d", X"d3", X"d9", X"c3", X"23", X"16", X"8e", X"f2", X"e1", X"51", X"f0", X"e8", X"40", X"75", X"12",
		X"30", X"0e", X"06", X"e1", X"c6", X"0f", X"ca", X"b8", X"fa", X"dc", X"1c", X"1e", X"1e", X"94", X"a9",
		X"d3", X"d9", X"6b", X"6e", X"8f", X"a3", X"5b", X"37", X"67", X"73", X"99", X"46", X"d7", X"47", X"0e",
		X"f7", X"ef", X"a7", X"b2", X"88", X"6c", X"a0", X"86", X"e2", X"13", X"22", X"3b", X"a4", X"8c", X"58",
		X"1f", X"99", X"4a", X"19", X"14", X"ed", X"60", X"46", X"ff", X"00", X"bb", X"f2", X"b2", X"b7", X"19",
		X"19", X"07", X"dc", X"b4", X"9f", X"8a", X"5f", X"19", X"fc", X"23", X"e1", X"8f", X"0c", X"6a", X"b3",
		X"69", X"d7", X"76", X"9a", X"35", X"95", X"c4", X"70", X"68", X"53", X"cb", X"a0", X"bc", X"16", X"f2",
		X"db", X"b2", X"cf", X"89", X"8c", X"b1", X"2a", X"34", X"db", X"d5", X"ae", X"42", X"e6", X"42", X"59",
		X"bc", X"d2", X"8a", X"5b", X"cc", X"6a", X"f1", X"ed", X"2a", X"ca", X"db", X"56", X"f0", X"37", X"89",
		X"7c", X"41", X"a9", X"c6", X"6e", X"b5", X"2f", X"ed", X"0b", X"34", X"37", X"52", X"b1", X"69", X"08",
		X"9a", X"57", X"32", X"fc", X"c4", X"e7", X"2c", X"46", X"49", X"eb", X"c9", X"f5", X"35", X"fa", X"f1",
		X"fb", X"2e", X"78", X"33", X"c2", X"9f", X"13", X"7f", X"64", X"af", X"87", X"3a", X"27", X"8e", X"f4",
		X"0b", X"3d", X"5f", X"4f", X"f8", X"85", X"15", X"fe", X"99", X"e2", X"3b", X"69", X"63", X"0b", X"1d",
		X"f4", X"36", X"52", X"5c", X"c3", X"68", X"db", X"53", X"02", X"29", X"a2", X"8e", X"de", X"dd", X"52",
		X"78", X"f6", X"ca", X"3c", X"88", X"8e", X"fc", X"c6", X"a4", X"70", X"50", X"9d", X"45", X"37", X"1a",
		X"4e", X"dd", X"1f", X"e0", X"d7", X"ae", X"b6", X"2a", X"14", X"d4", X"93", X"67", X"8b", X"7c", X"33",
		X"f8", X"bb", X"f0", X"3f", X"c4", X"bf", X"b3", X"de", X"8d", X"1f", X"8f", X"3c", X"4f", X"06", X"90",
		X"da", X"95", X"ee", X"ff", X"00", X"14", X"e9", X"ba", X"4e", X"9d", X"73", X"15", X"c6", X"9b", X"22",
		X"6a", X"29", X"9b", X"d9", X"ee", X"6d", X"22", X"4f", X"2e", X"3c", X"cb", X"04", X"d2", X"cb", X"88",
		X"f7", X"3c", X"fb", X"51", X"bc", X"c2", X"ae", X"9b", X"5a", X"bf", X"8d", X"3e", X"35", X"6b", X"3e",
		X"3f", X"f1", X"3e", X"b7", X"f0", X"e7", X"c4", X"5a", X"34", X"7a", X"4d", X"96", X"9b", X"6d", X"e2",
		X"1b", X"0d", X"52", X"47", X"7b", X"8d", X"3f", X"c4", X"17", X"82", X"26", X"68", X"ad", X"c4", X"f7",
		X"12", X"c7", X"6f", X"1c", X"2f", X"14", X"52", X"2c", X"d7", X"5e", X"63", X"15", X"f3", X"90", X"0c",
		X"6f", X"62", X"3c", X"07", X"f6", X"8f", X"f0", X"ae", X"8d", X"f0", X"43", X"5e", X"f1", X"85", X"9f",
		X"c2", X"a8", X"ee", X"fc", X"3b", X"0d", X"b7", X"c2", X"fd", X"2a", X"28", X"d6", X"da", X"fa", X"76",
		X"f9", X"35", X"0d", X"53", X"ec", X"97", X"aa", X"db", X"dd", X"b7", X"89", X"61", X"66", X"52", X"1b",
		X"38", X"63", X"bc", X"61", X"c0", X"6a", X"fa", X"4f", X"e0", X"35", X"85", X"be", X"8d", X"e0", X"2d",
		X"25", X"34", X"ff", X"00", X"35", X"21", X"b7", X"d3", X"7c", X"6f", X"61", X"15", X"bc", X"93", X"3c",
		X"b0", X"2c", X"1a", X"6e", X"bf", X"67", X"05", X"92", X"f9", X"4e", X"4a", X"66", X"38", X"de", X"41",
		X"bb", X"1b", X"98", X"bb", X"b3", X"96", X"66", X"24", X"fb", X"38", X"3a", X"8e", X"a5", X"47", X"2a",
		X"9b", X"ab", X"27", X"6e", X"ba", X"ff", X"00", X"c1", X"b9", X"4a", X"2d", X"fb", X"b7", X"d8", X"f9",
		X"cb", X"45", X"d6", X"fe", X"23", X"7c", X"24", X"f1", X"b7", X"8b", X"7e", X"28", X"7c", X"3d", X"f8",
		X"71", X"69", X"37", X"87", X"64", X"b0", X"d5", X"af", X"f4", X"6d", X"2a", X"eb", X"51", X"8a", X"58",
		X"f4", X"dd", X"08", X"24", X"91", X"a3", X"c3", X"e5", X"b1", X"77", X"8e", X"19", X"64", X"59", X"66",
		X"b6", X"8f", X"27", X"6d", X"bb", X"45", X"21", X"1e", X"5a", X"c8", X"bc", X"b7", X"ec", X"e7", X"f1",
		X"c3", X"c4", X"b6", X"9e", X"39", X"4f", X"16", X"fc", X"4b", X"8e", X"4d", X"6b", X"45", X"d5", X"64",
		X"6b", X"4b", X"61", X"2d", X"9d", X"b4", X"70", X"c7", X"2a", X"5c", X"5b", X"4c", X"d3", X"c4", X"1b",
		X"08", X"b2", X"a9", X"b5", X"85", X"9a", X"73", X"ca", X"3c", X"30", X"b1", X"93", X"78", X"dd", X"5f",
		X"a1", X"ba", X"bf", X"86", X"b4", X"2b", X"4f", X"8c", X"56", X"da", X"ad", X"be", X"9b", X"12", X"5c",
		X"e9", X"de", X"0d", X"d4", X"2d", X"6d", X"9b", X"92", X"ab", X"14", X"77", X"5a", X"64", X"88", X"85",
		X"4f", X"ca", X"c1", X"5d", X"98", X"8d", X"c0", X"e3", X"73", X"0e", X"84", X"8a", X"f8", X"03", X"fe",
		X"0a", X"0f", X"69", X"6b", X"63", X"fb", X"54", X"6a", X"90", X"58", X"c0", X"96", X"c9", X"a8", X"59",
		X"69", X"33", X"5c", X"88", X"46", X"cf", X"32", X"47", X"0f", X"0b", X"b1", X"c7", X"73", X"1c", X"31",
		X"a9", X"3d", X"4e", X"df", X"52", X"49", X"bc", X"6d", X"39", X"65", X"eb", X"da", X"d2", X"77", X"8a",
		X"96", X"cf", X"d3", X"ca", X"dd", X"cc", X"b9", X"a4", X"9d", X"ae", X"56", X"f1", X"2f", X"c4", X"2d",
		X"2f", X"5b", X"f0", X"dd", X"f7", X"89", X"a5", X"bc", X"36", X"de", X"22", X"d5", X"24", X"7d", X"43",
		X"52", X"98", X"ee", X"9e", X"df", X"4d", X"69", X"54", X"ec", X"58", X"d5", X"db", X"6a", X"dd", X"4a",
		X"c0", X"05", X"6e", X"91", X"a8", X"df", X"21", X"dd", X"b1", X"59", X"3e", X"1d", X"7c", X"7e", X"f8",
		X"a1", X"a3", X"f8", X"07", X"c3", X"7e", X"1f", X"f0", X"d4", X"5e", X"1a", X"b7", X"f0", X"7f", X"84",
		X"6f", X"ae", X"be", X"dd", X"1d", X"fc", X"b6", X"b6", X"f6", X"ba", X"a4", X"57", X"1b", X"d9", X"ac",
		X"24", X"86", X"77", X"df", X"75", X"0e", X"c9", X"6e", X"01", X"11", X"24", X"b2", X"37", X"da", X"30",
		X"e1", X"d9", X"93", X"77", X"85", X"f8", X"8f", X"52", X"d4", X"34", X"2d", X"5a", X"da", X"1d", X"1e",
		X"fa", X"e2", X"ce", X"38", X"d4", X"00", X"b0", X"c8", X"54", X"73", X"c9", X"27", X"d4", X"9c", X"9c",
		X"93", X"c9", X"ef", X"57", X"ee", X"2f", X"26", X"d7", X"74", X"3d", X"6b", X"52", X"d4", X"84", X"6f",
		X"75", X"61", X"30", X"48", X"25", X"8e", X"25", X"84", X"80", X"66", X"2a", X"77", X"6c", X"03", X"7f",
		X"03", X"f8", X"b3", X"dc", X"f5", X"26", X"be", X"52", X"38", X"ba", X"91", X"93", X"c4", X"c5", X"d9",
		X"cf", X"7b", X"69", X"be", X"bf", X"99", X"97", X"33", X"56", X"48", X"b5", X"e2", X"1b", X"9f", X"09",
		X"3d", X"ed", X"cd", X"8f", X"86", X"74", X"d3", X"a5", X"e8", X"e6", X"f1", X"ee", X"ed", X"ac", X"2d",
		X"e7", X"33", X"2d", X"b9", X"6e", X"06", X"e7", X"20", X"09", X"25", X"55", X"c2", X"b1", X"8c", X"79",
		X"65", X"95", X"ca", X"6e", X"52", X"09", X"f5", X"1b", X"1f", X"da", X"3f", X"c4", X"96", X"56", X"56",
		X"f6", X"76", X"ff", X"00", X"0d", X"b4", X"c6", X"8a", X"08", X"92", X"24", X"3b", X"e3", X"5c", X"aa",
		X"80", X"07", X"1b", X"b8", X"e0", X"74", X"ae", X"37", X"e2", X"2f", X"86", X"74", X"1d", X"1f", X"41",
		X"b4", X"9b", X"4c", X"d3", X"22", X"b7", X"70", X"96", X"e8", X"59", X"33", X"96", X"04", X"39", X"cb",
		X"73", X"f3", X"1c", X"a8", X"e4", X"e4", X"f5", X"e7", X"93", X"5e", X"cd", X"e1", X"8f", X"02", X"78",
		X"5a", X"f3", X"c3", X"7a", X"4d", X"dd", X"ce", X"9a", X"ef", X"34", X"f6", X"30", X"49", X"23", X"7d",
		X"a6", X"51", X"b9", X"9a", X"35", X"24", X"e0", X"36", X"3a", X"9a", X"f0", X"31", X"52", X"85", X"47",
		X"cd", X"35", X"7d", X"5e", X"f7", X"fd", X"19", X"dd", X"4a", X"b5", X"58", X"d4", X"92", X"52", X"3f",
		X"ff", X"d9"
	);

	-- Access 'stdout' model 'fifo_out'
	signal stdout_data : std_logic_vector(7 downto 0) := (others => '0');
	signal stdout_rdy : std_logic := '0';
	signal stdout_ack : std_logic := '0';
	signal stdout_vector_idx : natural := 0;
	signal stdout_vector : std_logic_vector(7 downto 0) := (others => '0');
	-- Test vectors
	constant stdout_vectors_nb : natural := 15932;
	type stdout_vec_type is array (0 to stdout_vectors_nb-1) of std_logic_vector(7 downto 0);
	constant stdout_vectors : stdout_vec_type := (
		X"bc", X"d1", X"be", X"99", X"8f", X"67", X"95", X"c0", X"ac", X"9d", X"bd", X"c0", X"a4", X"c3", X"bc",
		X"b5", X"c1", X"a7", X"bc", X"d2", X"b1", X"8e", X"25", X"0a", X"1f", X"28", X"27", X"34", X"20", X"1d",
		X"22", X"0e", X"0a", X"12", X"0e", X"1a", X"07", X"6c", X"b5", X"be", X"b5", X"7f", X"5b", X"63", X"49",
		X"24", X"0b", X"24", X"42", X"5d", X"5a", X"41", X"33", X"20", X"24", X"23", X"26", X"35", X"38", X"23",
		X"19", X"19", X"20", X"31", X"29", X"36", X"20", X"1f", X"1f", X"22", X"18", X"19", X"26", X"2b", X"20",
		X"0b", X"09", X"0d", X"14", X"19", X"17", X"11", X"10", X"12", X"1e", X"19", X"21", X"2d", X"24", X"1d",
		X"a6", X"c1", X"65", X"5a", X"aa", X"81", X"92", X"d5", X"a9", X"58", X"91", X"c7", X"cf", X"a5", X"89",
		X"71", X"c9", X"9b", X"8b", X"d1", X"bf", X"c9", X"ab", X"67", X"33", X"1d", X"11", X"09", X"1d", X"2b",
		X"21", X"24", X"18", X"0e", X"18", X"18", X"04", X"6c", X"b9", X"b4", X"ba", X"bc", X"b7", X"c3", X"c0",
		X"6c", X"30", X"4b", X"67", X"55", X"45", X"31", X"2e", X"37", X"2c", X"2a", X"32", X"33", X"29", X"1e",
		X"12", X"0e", X"1e", X"30", X"30", X"36", X"22", X"28", X"26", X"24", X"1f", X"1c", X"34", X"37", X"2d",
		X"0f", X"0e", X"10", X"17", X"15", X"0f", X"0b", X"11", X"19", X"1f", X"1a", X"2c", X"49", X"22", X"27",
		X"91", X"84", X"2e", X"b5", X"cd", X"d1", X"bb", X"aa", X"8c", X"38", X"34", X"8e", X"7a", X"b0", X"c6",
		X"53", X"9a", X"d7", X"c8", X"d1", X"b8", X"a4", X"c4", X"ae", X"80", X"37", X"59", X"4c", X"1c", X"26",
		X"2f", X"2e", X"23", X"1b", X"27", X"1f", X"10", X"3a", X"74", X"89", X"a9", X"b8", X"b4", X"af", X"a6",
		X"78", X"49", X"5b", X"61", X"54", X"20", X"24", X"3e", X"3a", X"28", X"29", X"30", X"2d", X"20", X"14",
		X"0f", X"10", X"0c", X"1b", X"18", X"24", X"28", X"10", X"22", X"18", X"16", X"21", X"3d", X"41", X"37",
		X"12", X"15", X"16", X"1d", X"13", X"12", X"0f", X"15", X"1c", X"21", X"1d", X"30", X"4b", X"24", X"26",
		X"6f", X"0f", X"3e", X"e2", X"cf", X"bb", X"cd", X"bc", X"3d", X"02", X"0d", X"1f", X"09", X"69", X"8c",
		X"31", X"18", X"bf", X"d1", X"c6", X"ba", X"b8", X"93", X"75", X"59", X"3a", X"8a", X"b3", X"87", X"3e",
		X"34", X"33", X"17", X"14", X"22", X"1c", X"1a", X"0a", X"2a", X"70", X"97", X"9d", X"8b", X"7a", X"71",
		X"36", X"4f", X"54", X"60", X"2e", X"13", X"20", X"35", X"3a", X"28", X"28", X"27", X"26", X"15", X"15",
		X"11", X"17", X"06", X"6e", X"65", X"0e", X"12", X"07", X"0f", X"1b", X"07", X"1b", X"40", X"46", X"3f",
		X"16", X"1e", X"20", X"26", X"16", X"08", X"0a", X"12", X"14", X"1a", X"1b", X"2b", X"3a", X"2c", X"28",
		X"8b", X"8c", X"81", X"9c", X"71", X"b1", X"d7", X"ae", X"6f", X"65", X"24", X"0e", X"14", X"8b", X"62",
		X"6a", X"51", X"25", X"61", X"df", X"c8", X"d9", X"95", X"99", X"94", X"83", X"46", X"92", X"b2", X"ac",
		X"83", X"50", X"0d", X"11", X"2b", X"10", X"12", X"14", X"18", X"62", X"82", X"a3", X"90", X"55", X"47",
		X"51", X"4e", X"58", X"44", X"1d", X"27", X"38", X"3b", X"31", X"28", X"29", X"27", X"14", X"0b", X"3f",
		X"50", X"01", X"59", X"b3", X"ba", X"60", X"00", X"25", X"0f", X"15", X"14", X"1b", X"40", X"4c", X"49",
		X"1d", X"1f", X"21", X"2b", X"22", X"0d", X"0c", X"13", X"10", X"10", X"0e", X"1c", X"26", X"3c", X"32",
		X"b3", X"c4", X"d9", X"84", X"37", X"79", X"d5", X"b4", X"b1", X"b7", X"ae", X"66", X"a1", X"b6", X"8c",
		X"93", X"c5", X"ce", X"a4", X"d6", X"d9", X"af", X"28", X"8d", X"ae", X"b7", X"7b", X"44", X"61", X"77",
		X"7b", X"7e", X"31", X"15", X"27", X"11", X"17", X"1c", X"0e", X"7b", X"95", X"c2", X"c1", X"5f", X"4b",
		X"49", X"46", X"3f", X"3b", X"32", X"30", X"37", X"3a", X"2a", X"30", X"36", X"20", X"24", X"0c", X"55",
		X"9f", X"6e", X"7d", X"b1", X"bb", X"89", X"19", X"36", X"3a", X"37", X"12", X"13", X"3b", X"4d", X"4c",
		X"22", X"1e", X"20", X"30", X"2f", X"22", X"12", X"0d", X"0d", X"0c", X"05", X"0c", X"12", X"34", X"39",
		X"88", X"86", X"af", X"d6", X"86", X"a1", X"be", X"8d", X"b1", X"bd", X"8d", X"a4", X"cb", X"b3", X"b9",
		X"90", X"49", X"8d", X"ce", X"94", X"b5", X"c0", X"71", X"45", X"95", X"b0", X"8d", X"74", X"53", X"2e",
		X"65", X"70", X"4f", X"1f", X"19", X"28", X"1e", X"1a", X"0c", X"62", X"a2", X"c3", X"d7", X"7a", X"37",
		X"41", X"3d", X"44", X"40", X"2e", X"44", X"41", X"43", X"50", X"38", X"24", X"2c", X"2f", X"1b", X"37",
		X"b1", X"c8", X"af", X"a9", X"b2", X"9c", X"72", X"7e", X"6b", X"3d", X"2e", X"32", X"3c", X"4e", X"4c",
		X"2e", X"2a", X"30", X"3b", X"3a", X"2d", X"19", X"14", X"16", X"1a", X"13", X"13", X"0f", X"38", X"3a",
		X"29", X"72", X"c4", X"c3", X"d0", X"c5", X"ba", X"b0", X"ae", X"cc", X"79", X"88", X"d0", X"cd", X"c9",
		X"56", X"0c", X"be", X"b4", X"b1", X"94", X"b2", X"dd", X"91", X"61", X"92", X"88", X"99", X"a9", X"8a",
		X"93", X"bf", X"a7", X"39", X"2f", X"a8", X"7c", X"21", X"05", X"36", X"bd", X"b4", X"c5", X"bc", X"88",
		X"44", X"36", X"3f", X"32", X"4e", X"53", X"4a", X"50", X"5a", X"3a", X"2c", X"3c", X"2d", X"2c", X"12",
		X"80", X"c2", X"b0", X"c9", X"cb", X"c4", X"af", X"8e", X"6b", X"3d", X"2c", X"3d", X"4a", X"56", X"53",
		X"3e", X"40", X"47", X"48", X"3f", X"3f", X"37", X"39", X"34", X"31", X"27", X"24", X"18", X"3d", X"39",
		X"13", X"4b", X"c2", X"a5", X"a8", X"ba", X"c4", X"bb", X"cb", X"cf", X"56", X"41", X"82", X"c0", X"d6",
		X"b8", X"90", X"ae", X"b4", X"d1", X"93", X"4c", X"6c", X"74", X"9b", X"9a", X"bb", X"ac", X"b3", X"b4",
		X"bb", X"c7", X"cc", X"39", X"36", X"a5", X"7f", X"2f", X"5a", X"43", X"bd", X"b3", X"aa", X"d6", X"c3",
		X"9f", X"67", X"28", X"20", X"40", X"61", X"42", X"35", X"35", X"43", X"4d", X"2e", X"2f", X"27", X"0a",
		X"35", X"7a", X"97", X"ca", X"d5", X"d6", X"bc", X"a1", X"91", X"6a", X"3c", X"3a", X"4e", X"5d", X"61",
		X"65", X"66", X"56", X"55", X"47", X"39", X"32", X"37", X"36", X"36", X"34", X"2b", X"28", X"15", X"16",
		X"71", X"0b", X"2e", X"42", X"68", X"8c", X"a4", X"a7", X"b1", X"d2", X"47", X"73", X"69", X"be", X"a3",
		X"b5", X"bb", X"b8", X"8e", X"b1", X"6b", X"cf", X"80", X"71", X"79", X"9c", X"99", X"8f", X"a1", X"9a",
		X"a5", X"b6", X"b6", X"37", X"2d", X"74", X"2a", X"34", X"78", X"5e", X"7d", X"b4", X"bb", X"ba", X"c7",
		X"bf", X"ba", X"4e", X"00", X"2b", X"60", X"76", X"52", X"13", X"4c", X"4c", X"47", X"37", X"1d", X"09",
		X"08", X"3b", X"6f", X"a8", X"bd", X"cd", X"bb", X"a6", X"8a", X"6f", X"32", X"29", X"37", X"4c", X"5e",
		X"6b", X"74", X"65", X"5c", X"48", X"33", X"32", X"2f", X"27", X"2b", X"25", X"1d", X"28", X"19", X"1b",
		X"64", X"44", X"33", X"2e", X"38", X"51", X"5c", X"98", X"b0", X"ca", X"47", X"8e", X"cf", X"c4", X"c5",
		X"90", X"b5", X"b5", X"69", X"78", X"4f", X"40", X"b3", X"70", X"66", X"61", X"40", X"3f", X"33", X"5e",
		X"b4", X"a4", X"93", X"25", X"44", X"a9", X"5e", X"64", X"61", X"8a", X"01", X"44", X"b2", X"b5", X"ad",
		X"a6", X"b6", X"a3", X"33", X"77", X"a5", X"bb", X"bb", X"41", X"27", X"4f", X"52", X"47", X"0f", X"0e",
		X"0a", X"0c", X"40", X"90", X"b9", X"b0", X"74", X"46", X"3c", X"29", X"27", X"19", X"17", X"2b", X"3f",
		X"56", X"6e", X"6e", X"64", X"4b", X"31", X"1b", X"20", X"1b", X"12", X"15", X"24", X"25", X"1d", X"20",
		X"5d", X"3e", X"22", X"1f", X"47", X"3e", X"66", X"af", X"90", X"6a", X"3a", X"c9", X"aa", X"bf", X"bd",
		X"a7", X"6e", X"aa", X"ae", X"86", X"79", X"54", X"a1", X"78", X"55", X"3e", X"40", X"2b", X"09", X"4e",
		X"ba", X"b9", X"aa", X"14", X"64", X"b4", X"9f", X"b0", X"ac", X"bd", X"64", X"6a", X"a9", X"aa", X"99",
		X"b4", X"bd", X"bb", X"bf", X"96", X"67", X"8a", X"9b", X"7d", X"31", X"4d", X"3d", X"3e", X"48", X"17",
		X"12", X"15", X"1b", X"27", X"52", X"50", X"35", X"35", X"47", X"54", X"3a", X"21", X"04", X"12", X"23",
		X"3f", X"65", X"78", X"6b", X"46", X"27", X"1c", X"1d", X"19", X"1c", X"18", X"20", X"21", X"22", X"1f",
		X"62", X"3b", X"20", X"11", X"22", X"1c", X"45", X"79", X"1a", X"2e", X"4c", X"ac", X"6b", X"13", X"8e",
		X"99", X"88", X"92", X"d6", X"a5", X"bb", X"cf", X"b3", X"7e", X"3f", X"51", X"26", X"2d", X"26", X"61",
		X"ad", X"b8", X"9b", X"18", X"64", X"ce", X"b0", X"c6", X"ce", X"e2", X"98", X"6b", X"81", X"99", X"92",
		X"bc", X"bb", X"aa", X"b3", X"b3", X"7c", X"9b", X"b3", X"9a", X"5d", X"49", X"41", X"51", X"42", X"39",
		X"14", X"3a", X"3c", X"24", X"2f", X"38", X"19", X"31", X"4a", X"5a", X"55", X"2c", X"08", X"0c", X"18",
		X"30", X"53", X"7a", X"78", X"57", X"25", X"1d", X"1c", X"17", X"17", X"14", X"1d", X"1f", X"17", X"14",
		X"61", X"33", X"09", X"0f", X"0e", X"10", X"17", X"58", X"20", X"25", X"4b", X"30", X"12", X"11", X"18",
		X"c5", X"c8", X"aa", X"c4", X"bf", X"ca", X"cd", X"b6", X"64", X"38", X"23", X"1c", X"71", X"5c", X"47",
		X"5d", X"56", X"56", X"22", X"4e", X"ba", X"c2", X"b6", X"c1", X"b4", X"a5", X"4e", X"56", X"7a", X"40",
		X"69", X"c3", X"a3", X"94", X"bc", X"94", X"96", X"96", X"76", X"78", X"5f", X"49", X"4d", X"4b", X"46",
		X"3f", X"4f", X"5f", X"40", X"52", X"3b", X"1f", X"14", X"2b", X"46", X"5d", X"54", X"1d", X"1d", X"2c",
		X"3e", X"4e", X"70", X"78", X"5d", X"2c", X"22", X"22", X"23", X"11", X"11", X"1c", X"14", X"17", X"1a",
		X"55", X"3a", X"15", X"18", X"1d", X"11", X"0d", X"1f", X"0d", X"15", X"59", X"1f", X"2d", X"13", X"15",
		X"92", X"e1", X"d2", X"ce", X"b9", X"42", X"a4", X"b7", X"bf", X"95", X"3c", X"42", X"77", X"34", X"4a",
		X"37", X"8e", X"9e", X"14", X"4b", X"9a", X"a1", X"c9", X"93", X"8a", X"b6", X"8f", X"7a", X"54", X"15",
		X"74", X"ae", X"ae", X"a8", X"c6", X"80", X"49", X"4e", X"a6", X"9f", X"4e", X"49", X"35", X"24", X"71",
		X"7c", X"58", X"80", X"7f", X"6a", X"42", X"09", X"17", X"14", X"29", X"4a", X"59", X"41", X"34", X"3e",
		X"49", X"3f", X"5b", X"6f", X"62", X"36", X"46", X"3d", X"3f", X"3c", X"32", X"1d", X"16", X"19", X"1c",
		X"25", X"50", X"19", X"17", X"10", X"04", X"0b", X"16", X"0d", X"16", X"56", X"1d", X"12", X"32", X"19",
		X"08", X"77", X"a3", X"a0", X"b9", X"a1", X"9e", X"bd", X"b3", X"84", X"77", X"74", X"27", X"81", X"ab",
		X"89", X"b4", X"ae", X"13", X"75", X"c2", X"c0", X"c1", X"ae", X"9f", X"77", X"a5", X"b1", X"a8", X"2c",
		X"79", X"a1", X"b9", X"c8", X"c2", X"a7", X"52", X"52", X"a2", X"a2", X"4a", X"33", X"37", X"0f", X"63",
		X"9c", X"76", X"7f", X"b1", X"a3", X"48", X"09", X"0d", X"0a", X"05", X"25", X"47", X"4d", X"46", X"6d",
		X"8d", X"7b", X"85", X"89", X"75", X"49", X"4f", X"45", X"53", X"50", X"52", X"43", X"2f", X"1c", X"1a",
		X"0d", X"4d", X"17", X"12", X"0f", X"10", X"10", X"22", X"21", X"15", X"55", X"0e", X"00", X"25", X"2c",
		X"00", X"b3", X"e1", X"bb", X"ce", X"d1", X"8d", X"95", X"4e", X"39", X"3f", X"48", X"81", X"9f", X"a4",
		X"6d", X"61", X"73", X"1f", X"24", X"5b", X"19", X"5d", X"d7", X"6c", X"64", X"b4", X"b5", X"78", X"44",
		X"52", X"a8", X"c3", X"c2", X"95", X"b9", X"b3", X"83", X"48", X"83", X"4b", X"37", X"2e", X"20", X"3d",
		X"90", X"96", X"81", X"c4", X"b6", X"79", X"57", X"51", X"06", X"05", X"14", X"26", X"38", X"64", X"99",
		X"ac", X"cc", X"cc", X"c6", X"d4", X"56", X"20", X"41", X"33", X"3b", X"39", X"3b", X"34", X"33", X"2c",
		X"2b", X"1e", X"20", X"14", X"32", X"46", X"31", X"13", X"1a", X"28", X"45", X"64", X"4b", X"32", X"28",
		X"12", X"64", X"c0", X"68", X"64", X"69", X"76", X"83", X"81", X"2a", X"4c", X"23", X"49", X"7c", X"92",
		X"68", X"01", X"1c", X"4b", X"62", X"c5", X"a6", X"b1", X"d4", X"c9", X"af", X"ae", X"c0", X"8e", X"63",
		X"21", X"57", X"d8", X"bd", X"c1", X"d1", X"b9", X"bc", X"7e", X"7e", X"5c", X"56", X"3a", X"23", X"1c",
		X"74", X"ae", X"b5", X"bc", X"b4", X"a6", X"88", X"56", X"10", X"01", X"00", X"06", X"17", X"3f", X"67",
		X"88", X"ae", X"c0", X"9b", X"c6", X"ad", X"23", X"10", X"2a", X"33", X"28", X"26", X"3a", X"2b", X"2c",
		X"1a", X"1d", X"19", X"0e", X"25", X"4b", X"23", X"3b", X"13", X"3b", X"3d", X"65", X"37", X"51", X"4f",
		X"1d", X"30", X"56", X"6d", X"51", X"42", X"bb", X"8f", X"b6", X"8e", X"0d", X"02", X"27", X"4e", X"90",
		X"69", X"1c", X"22", X"54", X"1b", X"5d", X"fd", X"a9", X"f2", X"5d", X"d8", X"a1", X"9b", X"c2", X"e7",
		X"8b", X"07", X"5b", X"cd", X"cc", X"e2", X"b8", X"df", X"ea", X"be", X"70", X"5c", X"2b", X"25", X"14",
		X"84", X"c2", X"c6", X"cb", X"ae", X"8a", X"3a", X"07", X"00", X"1a", X"66", X"6e", X"5b", X"79", X"78",
		X"84", X"6d", X"ab", X"a7", X"a5", X"d9", X"b0", X"52", X"4d", X"44", X"33", X"16", X"26", X"2c", X"2c",
		X"05", X"16", X"1d", X"1d", X"07", X"63", X"1e", X"8b", X"65", X"35", X"3c", X"64", X"87", X"4c", X"40",
		X"20", X"24", X"33", X"36", X"57", X"6f", X"93", X"f0", X"ba", X"ac", X"cd", X"2e", X"00", X"2e", X"15",
		X"0b", X"3e", X"25", X"2d", X"1a", X"00", X"2e", X"c2", X"ba", X"3c", X"ef", X"62", X"8c", X"c0", X"79",
		X"13", X"b2", X"a4", X"5e", X"b7", X"43", X"57", X"c2", X"c2", X"c4", X"be", X"53", X"22", X"20", X"38",
		X"55", X"ab", X"b6", X"af", X"ce", X"99", X"3d", X"01", X"06", X"40", X"a1", X"c6", X"b3", X"ac", X"b3",
		X"aa", X"70", X"a2", X"dd", X"bf", X"b9", X"b5", X"88", X"5a", X"56", X"39", X"1d", X"1b", X"2c", X"2b",
		X"35", X"14", X"0c", X"12", X"21", X"60", X"38", X"9c", X"8b", X"84", X"3d", X"2f", X"75", X"71", X"65",
		X"24", X"1b", X"05", X"3f", X"a6", X"7b", X"15", X"a3", X"cf", X"e0", X"b4", X"81", X"d4", X"9f", X"c1",
		X"cd", X"2a", X"14", X"33", X"17", X"1b", X"11", X"30", X"f0", X"34", X"b1", X"b1", X"95", X"40", X"01",
		X"8c", X"ba", X"b4", X"cc", X"d3", X"d5", X"65", X"bb", X"c6", X"96", X"3a", X"70", X"81", X"56", X"37",
		X"3f", X"4d", X"4a", X"66", X"92", X"9a", X"63", X"35", X"30", X"1c", X"57", X"b3", X"b1", X"af", X"b2",
		X"af", X"74", X"86", X"9d", X"b2", X"c1", X"b4", X"94", X"7d", X"55", X"1c", X"14", X"12", X"3a", X"3b",
		X"1f", X"2b", X"0a", X"47", X"b1", X"92", X"2d", X"99", X"76", X"b8", X"8d", X"33", X"1b", X"38", X"4d",
		X"2d", X"1e", X"48", X"91", X"9f", X"5a", X"58", X"a8", X"8e", X"b7", X"d4", X"56", X"ad", X"cc", X"c9",
		X"84", X"00", X"21", X"31", X"15", X"09", X"00", X"7d", X"be", X"3d", X"51", X"b1", X"5f", X"48", X"17",
		X"0f", X"60", X"ad", X"d6", X"b4", X"e5", X"da", X"ba", X"b9", X"df", X"48", X"92", X"a0", X"81", X"56",
		X"3e", X"4e", X"42", X"5d", X"6f", X"71", X"5a", X"49", X"52", X"4a", X"03", X"42", X"96", X"bf", X"b5",
		X"68", X"78", X"5a", X"74", X"72", X"7d", X"ab", X"7a", X"84", X"42", X"15", X"19", X"1b", X"3b", X"3c",
		X"25", X"21", X"0d", X"1a", X"c9", X"bf", X"34", X"aa", X"89", X"bd", X"d9", X"d0", X"98", X"1a", X"6f",
		X"28", X"0a", X"94", X"a9", X"a2", X"99", X"86", X"cc", X"cb", X"ab", X"92", X"3d", X"65", X"ca", X"8e",
		X"00", X"09", X"2c", X"36", X"13", X"0c", X"00", X"24", X"a7", X"52", X"1c", X"d9", X"7b", X"66", X"0c",
		X"35", X"17", X"00", X"2f", X"00", X"c3", X"c2", X"bc", X"ac", X"b0", X"ae", X"3d", X"65", X"9d", X"88",
		X"6d", X"28", X"2c", X"7d", X"92", X"93", X"80", X"4d", X"61", X"71", X"53", X"36", X"ac", X"be", X"a5",
		X"9f", X"bf", X"55", X"41", X"3f", X"21", X"2d", X"3f", X"3c", X"21", X"15", X"13", X"10", X"3f", X"3d",
		X"22", X"33", X"39", X"30", X"24", X"89", X"18", X"7a", X"5a", X"e6", X"c2", X"d2", X"be", X"50", X"2a",
		X"33", X"12", X"95", X"d3", X"9f", X"27", X"7b", X"ac", X"60", X"3f", X"09", X"4a", X"2a", X"94", X"e0",
		X"77", X"00", X"35", X"34", X"1e", X"00", X"2b", X"bd", X"75", X"5e", X"25", X"9f", X"9d", X"d6", X"67",
		X"16", X"1e", X"0d", X"3a", X"3c", X"2c", X"43", X"64", X"a8", X"a3", X"b3", X"36", X"8b", X"db", X"c1",
		X"71", X"44", X"8c", X"8f", X"8d", X"a5", X"79", X"7e", X"57", X"92", X"7c", X"5f", X"a6", X"a7", X"82",
		X"9c", X"bd", X"6c", X"2a", X"2b", X"29", X"11", X"28", X"1e", X"1d", X"17", X"13", X"12", X"3d", X"3c",
		X"0d", X"23", X"5e", X"7a", X"32", X"75", X"cd", X"ac", X"93", X"6c", X"dd", X"ba", X"b7", X"89", X"26",
		X"25", X"1f", X"6a", X"d0", X"9c", X"12", X"af", X"e5", X"8b", X"00", X"69", X"72", X"63", X"0c", X"92",
		X"8d", X"a2", X"34", X"2a", X"00", X"3e", X"b1", X"ba", X"88", X"5e", X"20", X"7b", X"92", X"d2", X"c1",
		X"6c", X"a8", X"91", X"08", X"c1", X"24", X"3d", X"45", X"3d", X"a6", X"9c", X"cb", X"7f", X"c3", X"e4",
		X"92", X"a9", X"8d", X"5a", X"88", X"6d", X"5f", X"62", X"5a", X"99", X"8f", X"56", X"52", X"61", X"60",
		X"63", X"7f", X"84", X"26", X"2e", X"24", X"1e", X"18", X"23", X"17", X"19", X"1b", X"0c", X"10", X"1e",
		X"0e", X"00", X"04", X"16", X"72", X"99", X"9e", X"ad", X"bc", X"bc", X"2f", X"70", X"f8", X"6d", X"cd",
		X"2e", X"22", X"4f", X"b5", X"6a", X"2c", X"b6", X"c9", X"8d", X"00", X"96", X"ac", X"7e", X"aa", X"a0",
		X"86", X"7a", X"6b", X"37", X"cc", X"6d", X"3e", X"98", X"eb", X"5c", X"26", X"86", X"65", X"b7", X"d9",
		X"94", X"98", X"9f", X"73", X"bf", X"b0", X"9b", X"90", X"5f", X"3e", X"34", X"ba", X"92", X"d8", X"b2",
		X"fb", X"60", X"49", X"7e", X"8a", X"38", X"61", X"37", X"67", X"78", X"7e", X"49", X"30", X"22", X"39",
		X"30", X"8d", X"8a", X"39", X"21", X"22", X"23", X"17", X"16", X"1f", X"1c", X"14", X"17", X"21", X"1e",
		X"2e", X"01", X"13", X"1d", X"1b", X"7c", X"a4", X"ac", X"ca", X"da", X"b0", X"64", X"18", X"6e", X"bd",
		X"32", X"2c", X"25", X"63", X"1d", X"1f", X"62", X"a4", X"30", X"47", X"c5", X"99", X"ca", X"a7", X"9c",
		X"c4", X"c0", X"38", X"80", X"d9", X"af", X"7d", X"99", X"31", X"6a", X"0f", X"80", X"ef", X"b6", X"c3",
		X"ab", X"5c", X"25", X"6e", X"56", X"76", X"94", X"62", X"37", X"22", X"1e", X"15", X"30", X"e8", X"d1",
		X"6a", X"57", X"6b", X"ac", X"1e", X"47", X"56", X"58", X"48", X"3e", X"31", X"42", X"2e", X"40", X"50",
		X"44", X"4c", X"6f", X"2d", X"2a", X"23", X"22", X"1c", X"1a", X"31", X"2b", X"16", X"1d", X"20", X"20",
		X"90", X"29", X"00", X"15", X"02", X"00", X"58", X"a0", X"a7", X"c0", X"a8", X"57", X"00", X"a9", X"eb",
		X"32", X"23", X"16", X"0c", X"62", X"00", X"17", X"3d", X"00", X"47", X"35", X"f0", X"90", X"ce", X"b2",
		X"bc", X"e1", X"c8", X"a7", X"ce", X"df", X"76", X"0c", X"4b", X"6d", X"24", X"51", X"e1", X"c2", X"90",
		X"b6", X"49", X"20", X"20", X"70", X"a7", X"5d", X"32", X"2c", X"1e", X"11", X"33", X"2b", X"5d", X"75",
		X"71", X"49", X"d2", X"a2", X"63", X"57", X"57", X"41", X"22", X"22", X"16", X"15", X"23", X"48", X"67",
		X"63", X"3a", X"38", X"2f", X"2d", X"28", X"1a", X"1e", X"22", X"3e", X"39", X"20", X"25", X"1e", X"1e",
		X"b7", X"70", X"00", X"08", X"0b", X"1a", X"00", X"77", X"cd", X"94", X"d2", X"00", X"3c", X"e1", X"53",
		X"3a", X"23", X"1e", X"06", X"25", X"3d", X"07", X"69", X"1f", X"24", X"07", X"59", X"e5", X"ab", X"ac",
		X"c3", X"db", X"d3", X"af", X"b1", X"db", X"90", X"4a", X"2f", X"6a", X"25", X"32", X"c2", X"bc", X"64",
		X"53", X"19", X"40", X"31", X"bb", X"af", X"84", X"19", X"2b", X"19", X"20", X"30", X"1e", X"4a", X"6c",
		X"5a", X"8b", X"d2", X"c5", X"83", X"6a", X"4f", X"2a", X"56", X"40", X"23", X"24", X"26", X"44", X"5d",
		X"57", X"67", X"36", X"57", X"29", X"29", X"15", X"18", X"1d", X"3d", X"3a", X"26", X"37", X"14", X"1e",
		X"91", X"4c", X"05", X"0a", X"02", X"23", X"00", X"91", X"bf", X"d7", X"3b", X"05", X"96", X"b3", X"89",
		X"2e", X"2c", X"18", X"09", X"18", X"46", X"3e", X"15", X"0b", X"41", X"8d", X"57", X"7f", X"ad", X"8b",
		X"a9", X"6c", X"d4", X"b5", X"96", X"c2", X"ca", X"9a", X"52", X"3a", X"50", X"3c", X"59", X"8d", X"54",
		X"00", X"68", X"68", X"1a", X"52", X"a1", X"55", X"0c", X"10", X"3c", X"4c", X"48", X"02", X"52", X"7c",
		X"61", X"a2", X"f1", X"b9", X"74", X"91", X"2a", X"31", X"58", X"44", X"2a", X"14", X"1b", X"41", X"55",
		X"64", X"4f", X"5d", X"3a", X"4c", X"1e", X"16", X"15", X"1c", X"3d", X"3a", X"25", X"41", X"20", X"1c",
		X"63", X"28", X"05", X"09", X"0b", X"17", X"2a", X"dc", X"c4", X"ff", X"00", X"1a", X"e2", X"a4", X"82",
		X"6e", X"1d", X"1f", X"00", X"1f", X"46", X"29", X"25", X"27", X"66", X"7e", X"9c", X"d1", X"9e", X"d7",
		X"f9", X"e2", X"de", X"c3", X"e8", X"e2", X"ca", X"a3", X"5d", X"3f", X"54", X"33", X"83", X"9d", X"00",
		X"8b", X"4b", X"72", X"3b", X"0b", X"7c", X"5e", X"1c", X"45", X"6e", X"61", X"2f", X"2c", X"91", X"68",
		X"63", X"27", X"b5", X"bc", X"b9", X"b7", X"36", X"12", X"27", X"2e", X"43", X"2d", X"07", X"67", X"a3",
		X"86", X"6d", X"4d", X"4b", X"28", X"1a", X"16", X"18", X"23", X"3e", X"40", X"25", X"32", X"20", X"1f",
		X"87", X"68", X"0a", X"02", X"14", X"14", X"1a", X"00", X"1e", X"0e", X"15", X"4f", X"88", X"6c", X"65",
		X"26", X"38", X"16", X"19", X"1f", X"41", X"3d", X"0e", X"16", X"3b", X"77", X"3a", X"52", X"62", X"4a",
		X"29", X"9d", X"c8", X"48", X"52", X"da", X"9d", X"a6", X"79", X"52", X"71", X"11", X"9e", X"d1", X"92",
		X"7f", X"3e", X"7e", X"38", X"07", X"46", X"62", X"61", X"49", X"49", X"62", X"04", X"a6", X"6a", X"75",
		X"2a", X"25", X"01", X"b6", X"cb", X"b2", X"3c", X"1e", X"19", X"2d", X"37", X"29", X"16", X"40", X"b7",
		X"c5", X"b4", X"61", X"42", X"27", X"22", X"15", X"16", X"28", X"38", X"44", X"2c", X"1f", X"1f", X"21",
		X"55", X"20", X"3e", X"00", X"14", X"11", X"23", X"2c", X"13", X"17", X"00", X"93", X"d0", X"49", X"55",
		X"0e", X"46", X"09", X"24", X"25", X"3a", X"4e", X"17", X"2f", X"04", X"0b", X"14", X"03", X"3e", X"41",
		X"12", X"92", X"c5", X"86", X"6f", X"c0", X"df", X"ba", X"a0", X"7f", X"7d", X"3c", X"ab", X"d2", X"d4",
		X"cf", X"a8", X"ae", X"90", X"bf", X"00", X"94", X"78", X"23", X"42", X"1d", X"4f", X"b6", X"5f", X"47",
		X"19", X"5e", X"72", X"47", X"a6", X"bf", X"93", X"60", X"18", X"14", X"2f", X"1f", X"27", X"28", X"70",
		X"a8", X"d1", X"98", X"4d", X"27", X"11", X"0c", X"1d", X"33", X"41", X"4a", X"2c", X"0f", X"07", X"15",
		X"51", X"42", X"0c", X"28", X"00", X"0d", X"5a", X"18", X"13", X"23", X"01", X"95", X"2f", X"5c", X"5b",
		X"07", X"44", X"0a", X"2c", X"1c", X"1c", X"5f", X"00", X"a0", X"6a", X"0e", X"1d", X"0c", X"45", X"2b",
		X"15", X"f5", X"bf", X"7a", X"c3", X"e5", X"d1", X"cf", X"9b", X"61", X"8a", X"fe", X"af", X"76", X"f7",
		X"d9", X"d9", X"b7", X"5e", X"6b", X"73", X"42", X"66", X"8a", X"0d", X"10", X"9c", X"80", X"2f", X"16",
		X"0f", X"2c", X"a2", X"8a", X"9b", X"a5", X"a7", X"ac", X"58", X"03", X"23", X"1f", X"87", X"86", X"b4",
		X"9b", X"c0", X"be", X"a5", X"35", X"09", X"11", X"1c", X"35", X"4b", X"4e", X"46", X"37", X"1e", X"26",
		X"39", X"71", X"07", X"21", X"0a", X"1f", X"45", X"17", X"2a", X"0d", X"1c", X"08", X"01", X"37", X"1b",
		X"3b", X"3d", X"1b", X"29", X"21", X"0d", X"25", X"28", X"84", X"8f", X"08", X"16", X"10", X"2c", X"58",
		X"54", X"48", X"98", X"a8", X"ac", X"c1", X"93", X"c9", X"b2", X"65", X"00", X"e0", X"e7", X"fa", X"30",
		X"03", X"c1", X"e9", X"3c", X"4e", X"21", X"9f", X"8f", X"d4", X"00", X"32", X"00", X"09", X"0b", X"4b",
		X"27", X"41", X"43", X"c6", X"c8", X"91", X"38", X"52", X"4f", X"14", X"32", X"53", X"27", X"69", X"33",
		X"46", X"b9", X"d2", X"d0", X"bd", X"39", X"0f", X"19", X"29", X"3b", X"48", X"50", X"70", X"1f", X"24",
		X"40", X"72", X"61", X"00", X"18", X"58", X"95", X"1c", X"0f", X"2e", X"10", X"09", X"36", X"3e", X"01",
		X"00", X"6e", X"3f", X"10", X"1b", X"21", X"38", X"17", X"11", X"00", X"2b", X"2e", X"42", X"3e", X"0c",
		X"7f", X"a7", X"bd", X"39", X"fb", X"e3", X"7a", X"02", X"00", X"07", X"44", X"36", X"5f", X"50", X"f7",
		X"a5", X"d4", X"40", X"6f", X"3e", X"db", X"32", X"7f", X"2b", X"53", X"38", X"24", X"11", X"31", X"42",
		X"7b", X"6f", X"79", X"91", X"7f", X"af", X"bb", X"54", X"60", X"5f", X"0f", X"21", X"38", X"82", X"82",
		X"ce", X"a8", X"bb", X"ce", X"b3", X"90", X"2d", X"2b", X"1b", X"18", X"4b", X"6e", X"7a", X"23", X"1d",
		X"5e", X"49", X"4b", X"86", X"0d", X"22", X"50", X"4a", X"0b", X"79", X"6f", X"2d", X"33", X"1d", X"22",
		X"be", X"d5", X"7a", X"11", X"19", X"19", X"0b", X"6e", X"73", X"21", X"2c", X"42", X"0a", X"2b", X"05",
		X"42", X"73", X"85", X"39", X"4a", X"f4", X"82", X"00", X"23", X"10", X"14", X"59", X"2a", X"3c", X"e6",
		X"db", X"4e", X"c5", X"eb", X"8b", X"93", X"2e", X"0a", X"7a", X"75", X"6f", X"5a", X"36", X"38", X"43",
		X"52", X"3a", X"10", X"8b", X"91", X"9e", X"d2", X"67", X"12", X"25", X"30", X"23", X"20", X"25", X"09",
		X"21", X"23", X"78", X"a1", X"af", X"79", X"44", X"2e", X"0e", X"16", X"38", X"67", X"7a", X"47", X"5c",
		X"57", X"53", X"00", X"5c", X"7f", X"14", X"2c", X"0f", X"76", X"7c", X"79", X"50", X"2f", X"53", X"95",
		X"8c", X"b6", X"41", X"11", X"1a", X"31", X"41", X"66", X"ba", X"74", X"16", X"82", X"0d", X"00", X"3f",
		X"28", X"37", X"18", X"65", X"0a", X"1c", X"82", X"02", X"15", X"2e", X"08", X"2f", X"3a", X"7a", X"fb",
		X"13", X"6a", X"d0", X"b4", X"d4", X"65", X"06", X"37", X"5c", X"3e", X"7d", X"41", X"59", X"27", X"22",
		X"1e", X"02", X"21", X"6f", X"56", X"77", X"d5", X"00", X"a3", X"5d", X"11", X"19", X"23", X"1b", X"1b",
		X"25", X"23", X"3f", X"69", X"aa", X"7d", X"32", X"18", X"02", X"10", X"2b", X"52", X"4e", X"62", X"61",
		X"58", X"12", X"1b", X"00", X"6f", X"7c", X"17", X"22", X"8f", X"d7", X"9c", X"b9", X"9f", X"7c", X"6e",
		X"5c", X"a1", X"40", X"16", X"0f", X"3b", X"42", X"41", X"4e", X"39", X"23", X"16", X"2a", X"0c", X"58",
		X"00", X"17", X"21", X"77", X"53", X"2b", X"00", X"12", X"20", X"36", X"16", X"32", X"37", X"03", X"25",
		X"9d", X"40", X"00", X"0b", X"92", X"16", X"42", X"63", X"44", X"5c", X"4e", X"46", X"a7", X"1a", X"18",
		X"07", X"0c", X"2c", X"3c", X"05", X"57", X"90", X"34", X"c2", X"aa", X"55", X"19", X"1c", X"1e", X"0f",
		X"19", X"16", X"15", X"35", X"7c", X"7e", X"52", X"36", X"0c", X"1c", X"24", X"38", X"3d", X"67", X"6b",
		X"87", X"0d", X"19", X"29", X"18", X"8e", X"2d", X"1c", X"13", X"f3", X"ca", X"ba", X"aa", X"eb", X"60",
		X"6f", X"8c", X"50", X"2c", X"08", X"23", X"15", X"64", X"14", X"0f", X"09", X"00", X"0b", X"25", X"00",
		X"1f", X"01", X"67", X"8e", X"64", X"00", X"0c", X"56", X"28", X"68", X"3e", X"0c", X"14", X"30", X"32",
		X"33", X"13", X"35", X"8e", X"13", X"3c", X"54", X"64", X"43", X"3f", X"5d", X"58", X"02", X"29", X"16",
		X"16", X"1c", X"2a", X"32", X"28", X"2c", X"23", X"56", X"78", X"8b", X"77", X"39", X"12", X"14", X"08",
		X"02", X"12", X"16", X"07", X"26", X"33", X"43", X"3a", X"3c", X"5b", X"26", X"30", X"47", X"6a", X"72",
		X"a8", X"f8", X"46", X"14", X"29", X"00", X"13", X"38", X"6d", X"30", X"d1", X"bd", X"9c", X"79", X"fb",
		X"ac", X"ca", X"75", X"82", X"73", X"3e", X"11", X"51", X"10", X"2b", X"bf", X"a5", X"43", X"02", X"12",
		X"30", X"b2", X"a0", X"72", X"00", X"8f", X"cc", X"bb", X"a9", X"2b", X"28", X"24", X"2e", X"23", X"4e",
		X"39", X"06", X"11", X"56", X"b4", X"1e", X"67", X"1c", X"17", X"73", X"62", X"3e", X"14", X"41", X"3a",
		X"37", X"48", X"56", X"52", X"51", X"50", X"41", X"17", X"39", X"5c", X"9a", X"40", X"61", X"4e", X"3a",
		X"28", X"21", X"2b", X"5b", X"27", X"19", X"0a", X"20", X"49", X"48", X"21", X"31", X"38", X"0c", X"00",
		X"4e", X"8c", X"be", X"00", X"5c", X"6c", X"12", X"0d", X"8b", X"c4", X"c7", X"d7", X"3a", X"4a", X"5d",
		X"d7", X"ad", X"60", X"3a", X"55", X"5f", X"15", X"31", X"52", X"00", X"66", X"db", X"be", X"96", X"03",
		X"97", X"7f", X"9e", X"9d", X"00", X"cd", X"dd", X"ad", X"bc", X"67", X"2b", X"30", X"24", X"48", X"5b",
		X"7b", X"6b", X"38", X"09", X"5d", X"02", X"58", X"0e", X"51", X"60", X"49", X"3c", X"14", X"3e", X"2d",
		X"36", X"44", X"29", X"39", X"1f", X"18", X"3c", X"5a", X"08", X"34", X"53", X"81", X"c3", X"81", X"5d",
		X"4e", X"58", X"83", X"6c", X"68", X"34", X"1d", X"2f", X"59", X"4d", X"33", X"34", X"54", X"01", X"03",
		X"5a", X"46", X"82", X"01", X"8a", X"c1", X"cc", X"85", X"9f", X"af", X"b8", X"dc", X"4d", X"67", X"b6",
		X"b9", X"d1", X"83", X"68", X"2c", X"30", X"2d", X"1a", X"4a", X"16", X"00", X"88", X"df", X"bb", X"b4",
		X"a2", X"44", X"e2", X"39", X"31", X"a9", X"98", X"d6", X"d6", X"b2", X"15", X"32", X"2c", X"3c", X"35",
		X"51", X"67", X"3d", X"26", X"20", X"16", X"32", X"02", X"43", X"ac", X"b7", X"b1", X"1b", X"23", X"17",
		X"0f", X"0e", X"72", X"50", X"28", X"2d", X"1c", X"0c", X"09", X"56", X"ac", X"af", X"b7", X"b7", X"7d",
		X"57", X"7d", X"58", X"82", X"5a", X"3b", X"12", X"41", X"6f", X"4e", X"25", X"22", X"3c", X"01", X"05",
		X"0c", X"1e", X"08", X"11", X"17", X"7c", X"c4", X"df", X"d4", X"92", X"79", X"c6", X"e6", X"e6", X"a2",
		X"d4", X"83", X"43", X"23", X"27", X"0e", X"1e", X"11", X"26", X"2b", X"ba", X"c0", X"b3", X"da", X"b8",
		X"d8", X"f9", X"1e", X"16", X"05", X"2b", X"ad", X"a5", X"9c", X"00", X"35", X"05", X"3a", X"34", X"44",
		X"67", X"1f", X"29", X"0e", X"10", X"50", X"20", X"0e", X"63", X"f8", X"c3", X"56", X"68", X"bc", X"ca",
		X"57", X"52", X"b6", X"8c", X"59", X"14", X"12", X"12", X"2f", X"30", X"6c", X"e1", X"b0", X"c6", X"ce",
		X"62", X"61", X"75", X"5a", X"47", X"29", X"0e", X"2a", X"63", X"35", X"1d", X"1c", X"29", X"07", X"00",
		X"1f", X"66", X"1a", X"36", X"09", X"00", X"9c", X"c5", X"e3", X"c7", X"cb", X"c8", X"eb", X"c2", X"8a",
		X"ca", X"9f", X"0e", X"2f", X"20", X"00", X"34", X"24", X"0c", X"6c", X"96", X"a4", X"b3", X"b3", X"62",
		X"9d", X"cf", X"01", X"0e", X"00", X"67", X"76", X"98", X"9f", X"00", X"22", X"99", X"60", X"4d", X"7f",
		X"12", X"04", X"67", X"13", X"1a", X"4e", X"40", X"a1", X"e5", X"34", X"00", X"00", X"44", X"a9", X"82",
		X"e7", X"48", X"d0", X"c5", X"7c", X"05", X"2e", X"5d", X"2f", X"47", X"54", X"37", X"e5", X"ca", X"cc",
		X"61", X"71", X"96", X"9a", X"88", X"8a", X"84", X"7d", X"34", X"49", X"16", X"4b", X"29", X"16", X"00",
		X"59", X"4b", X"38", X"49", X"4c", X"88", X"71", X"e2", X"b5", X"86", X"b0", X"d6", X"d6", X"67", X"96",
		X"87", X"d5", X"00", X"2f", X"12", X"05", X"0f", X"35", X"18", X"1c", X"3f", X"7f", X"c6", X"c5", X"ab",
		X"a1", X"db", X"cc", X"1e", X"00", X"75", X"5d", X"6e", X"9a", X"34", X"95", X"5e", X"67", X"8f", X"91",
		X"00", X"7f", X"92", X"7d", X"43", X"b3", X"b4", X"6b", X"00", X"09", X"59", X"c3", X"00", X"d1", X"9a",
		X"8c", X"c3", X"97", X"eb", X"a9", X"02", X"2d", X"31", X"47", X"9a", X"94", X"b0", X"bd", X"da", X"6b",
		X"47", X"bc", X"c7", X"97", X"4b", X"35", X"50", X"4a", X"32", X"44", X"15", X"44", X"38", X"04", X"0b",
		X"20", X"21", X"4d", X"87", X"c5", X"c0", X"b4", X"93", X"cf", X"5b", X"93", X"8d", X"c3", X"b6", X"61",
		X"64", X"93", X"01", X"2c", X"14", X"0c", X"0d", X"08", X"21", X"20", X"19", X"1e", X"52", X"73", X"96",
		X"d2", X"c0", X"df", X"d6", X"00", X"2d", X"c6", X"b1", X"b9", X"dc", X"57", X"5c", X"84", X"34", X"a9",
		X"ba", X"9a", X"a6", X"3a", X"29", X"58", X"2d", X"14", X"18", X"57", X"ff", X"52", X"a2", X"be", X"e6",
		X"d4", X"c0", X"c1", X"f1", X"53", X"13", X"2e", X"3e", X"81", X"b4", X"a8", X"b6", X"e4", X"ed", X"65",
		X"07", X"ae", X"bf", X"ab", X"a4", X"6d", X"43", X"0a", X"3b", X"3c", X"1b", X"1f", X"36", X"0f", X"0c",
		X"55", X"1f", X"89", X"5c", X"ad", X"ca", X"c0", X"bc", X"eb", X"1a", X"5b", X"dd", X"9f", X"d0", X"b5",
		X"18", X"0b", X"13", X"0c", X"12", X"04", X"0e", X"41", X"19", X"28", X"1a", X"6e", X"4c", X"86", X"6d",
		X"cb", X"c0", X"a0", X"ab", X"43", X"00", X"f7", X"c7", X"d4", X"f1", X"a6", X"8d", X"8d", X"4a", X"1c",
		X"d9", X"ce", X"bf", X"0b", X"40", X"30", X"67", X"64", X"3c", X"3c", X"e6", X"7b", X"31", X"83", X"7a",
		X"ae", X"d7", X"00", X"77", X"68", X"00", X"6b", X"88", X"57", X"5c", X"74", X"82", X"4f", X"62", X"f9",
		X"82", X"cf", X"d5", X"a0", X"00", X"00", X"13", X"21", X"3a", X"4d", X"29", X"27", X"3f", X"11", X"12",
		X"57", X"48", X"78", X"59", X"4a", X"de", X"dd", X"af", X"b6", X"d3", X"df", X"ab", X"e1", X"c1", X"88",
		X"08", X"0c", X"0b", X"0f", X"00", X"0d", X"01", X"52", X"19", X"22", X"2d", X"af", X"50", X"9b", X"3e",
		X"a3", X"a2", X"85", X"00", X"8d", X"ac", X"c0", X"c8", X"47", X"92", X"f8", X"c3", X"8c", X"b5", X"f0",
		X"9d", X"d8", X"d3", X"02", X"55", X"71", X"59", X"1a", X"a0", X"e0", X"a8", X"99", X"61", X"51", X"c1",
		X"2a", X"c9", X"03", X"d1", X"be", X"5a", X"47", X"81", X"59", X"3f", X"3f", X"6a", X"04", X"04", X"d2",
		X"b1", X"d6", X"9c", X"ec", X"26", X"0b", X"07", X"19", X"5f", X"60", X"29", X"31", X"3d", X"40", X"81",
		X"36", X"7c", X"67", X"60", X"5f", X"b9", X"12", X"93", X"d0", X"b8", X"a0", X"b9", X"a8", X"d1", X"00",
		X"0f", X"16", X"07", X"15", X"1a", X"1b", X"15", X"04", X"1e", X"18", X"8d", X"a5", X"bc", X"6d", X"2d",
		X"7e", X"79", X"8f", X"b4", X"ba", X"c1", X"e7", X"a4", X"44", X"08", X"a4", X"c1", X"71", X"7c", X"8d",
		X"af", X"a8", X"e3", X"7e", X"24", X"34", X"00", X"a0", X"88", X"bb", X"cb", X"6a", X"aa", X"52", X"3b",
		X"38", X"cb", X"e8", X"aa", X"98", X"62", X"2a", X"2c", X"4f", X"62", X"84", X"39", X"0b", X"58", X"c6",
		X"c1", X"ad", X"56", X"a5", X"f6", X"3f", X"21", X"0c", X"49", X"38", X"2a", X"29", X"31", X"7a", X"7c",
		X"6d", X"69", X"51", X"54", X"16", X"48", X"41", X"94", X"c3", X"dc", X"b8", X"d3", X"87", X"ca", X"34",
		X"00", X"0e", X"20", X"2e", X"2f", X"2c", X"19", X"23", X"1d", X"19", X"26", X"44", X"08", X"39", X"4e",
		X"59", X"87", X"2c", X"8b", X"a5", X"be", X"aa", X"ca", X"59", X"c7", X"c1", X"c8", X"88", X"80", X"9b",
		X"62", X"24", X"c5", X"ea", X"3a", X"00", X"25", X"48", X"72", X"ef", X"a1", X"35", X"00", X"13", X"00",
		X"3f", X"a3", X"9a", X"b8", X"96", X"59", X"62", X"68", X"66", X"7b", X"4a", X"07", X"59", X"06", X"7e",
		X"e8", X"38", X"11", X"3e", X"c6", X"75", X"69", X"43", X"25", X"1c", X"2b", X"32", X"1c", X"83", X"8d",
		X"2f", X"1c", X"23", X"5b", X"46", X"23", X"10", X"16", X"ce", X"bc", X"41", X"54", X"c8", X"8e", X"6d",
		X"1a", X"25", X"15", X"06", X"1d", X"05", X"1e", X"0f", X"11", X"1f", X"0b", X"0b", X"2b", X"3e", X"26",
		X"08", X"14", X"5e", X"66", X"b2", X"a1", X"9c", X"92", X"eb", X"ad", X"9d", X"87", X"6f", X"62", X"18",
		X"27", X"23", X"26", X"d4", X"73", X"00", X"30", X"3f", X"14", X"ee", X"00", X"05", X"0c", X"01", X"12",
		X"22", X"86", X"8f", X"cf", X"3e", X"55", X"61", X"7d", X"9a", X"40", X"00", X"34", X"09", X"23", X"3a",
		X"64", X"16", X"13", X"19", X"66", X"d6", X"31", X"2e", X"20", X"37", X"34", X"2e", X"31", X"8c", X"89",
		X"3b", X"17", X"08", X"57", X"6e", X"00", X"17", X"02", X"1a", X"a2", X"25", X"59", X"31", X"be", X"76",
		X"4f", X"03", X"0b", X"11", X"15", X"15", X"0b", X"15", X"04", X"2e", X"11", X"17", X"2d", X"33", X"2e",
		X"1a", X"36", X"00", X"0d", X"fe", X"e9", X"b8", X"d0", X"96", X"f0", X"a8", X"90", X"53", X"08", X"04",
		X"ec", X"cc", X"06", X"b8", X"00", X"22", X"3b", X"34", X"0f", X"00", X"19", X"2d", X"03", X"0b", X"37",
		X"1c", X"68", X"76", X"b6", X"1b", X"44", X"5e", X"9e", X"82", X"0a", X"76", X"3b", X"1e", X"29", X"3f",
		X"15", X"12", X"2b", X"2c", X"0b", X"60", X"07", X"2c", X"33", X"33", X"2d", X"33", X"35", X"6d", X"93",
		X"44", X"00", X"01", X"00", X"5b", X"41", X"07", X"0a", X"4b", X"6f", X"4a", X"18", X"c7", X"8f", X"8d",
		X"63", X"00", X"0a", X"2f", X"0c", X"16", X"19", X"10", X"10", X"26", X"0a", X"05", X"3c", X"59", X"08",
		X"15", X"44", X"12", X"37", X"eb", X"db", X"ff", X"c3", X"6b", X"ff", X"d3", X"c0", X"7a", X"0b", X"a3",
		X"a6", X"b2", X"17", X"4c", X"23", X"21", X"4f", X"19", X"30", X"0e", X"2c", X"0d", X"0d", X"13", X"07",
		X"1a", X"3c", X"47", X"53", X"1b", X"33", X"85", X"7b", X"00", X"5d", X"68", X"13", X"27", X"20", X"20",
		X"1f", X"00", X"02", X"15", X"68", X"06", X"8c", X"2b", X"23", X"20", X"2a", X"21", X"36", X"88", X"90",
		X"13", X"18", X"06", X"00", X"02", X"2f", X"04", X"13", X"45", X"58", X"62", X"84", X"db", X"c7", X"61",
		X"74", X"53", X"00", X"12", X"12", X"08", X"14", X"1b", X"0c", X"0e", X"0d", X"14", X"43", X"04", X"0c",
		X"2f", X"09", X"19", X"10", X"4c", X"ac", X"55", X"17", X"19", X"62", X"c4", X"b8", X"4a", X"13", X"b1",
		X"8d", X"da", X"f2", X"5b", X"bb", X"80", X"55", X"6b", X"d8", X"5c", X"00", X"10", X"0f", X"0b", X"39",
		X"55", X"12", X"35", X"92", X"17", X"56", X"55", X"03", X"58", X"3a", X"20", X"33", X"1d", X"10", X"0a",
		X"2a", X"c8", X"9b", X"a8", X"24", X"61", X"15", X"16", X"1b", X"1d", X"31", X"2a", X"1d", X"98", X"9d",
		X"1a", X"0b", X"0f", X"0a", X"0c", X"0c", X"0a", X"19", X"50", X"50", X"4d", X"1b", X"5f", X"a1", X"73",
		X"68", X"15", X"11", X"0c", X"0f", X"28", X"0e", X"12", X"0d", X"04", X"73", X"d4", X"6d", X"c0", X"21",
		X"1e", X"37", X"2e", X"1b", X"0f", X"4f", X"20", X"de", X"3e", X"08", X"06", X"8f", X"a8", X"a0", X"ac",
		X"b2", X"b3", X"55", X"55", X"41", X"cd", X"78", X"37", X"89", X"d1", X"0b", X"0e", X"00", X"4d", X"78",
		X"22", X"27", X"4b", X"31", X"29", X"34", X"12", X"2b", X"5b", X"43", X"0e", X"0f", X"06", X"16", X"1a",
		X"6b", X"3f", X"1c", X"00", X"27", X"20", X"18", X"1d", X"14", X"20", X"1f", X"27", X"2d", X"98", X"9b",
		X"0f", X"0d", X"00", X"00", X"0e", X"0c", X"04", X"22", X"3e", X"35", X"5d", X"38", X"49", X"06", X"27",
		X"78", X"6e", X"00", X"10", X"00", X"00", X"09", X"0d", X"00", X"20", X"bc", X"28", X"cf", X"f3", X"e2",
		X"00", X"06", X"0e", X"14", X"60", X"2f", X"18", X"b3", X"f8", X"2b", X"06", X"56", X"dc", X"96", X"b3",
		X"cf", X"a3", X"a2", X"8a", X"cc", X"d2", X"4a", X"2b", X"c6", X"a6", X"be", X"d3", X"ae", X"07", X"34",
		X"27", X"22", X"38", X"1e", X"1f", X"0b", X"33", X"3f", X"37", X"3b", X"57", X"53", X"46", X"2c", X"32",
		X"1b", X"20", X"22", X"23", X"20", X"26", X"1f", X"21", X"1a", X"3b", X"39", X"2d", X"34", X"43", X"49",
		X"00", X"00", X"06", X"03", X"0b", X"08", X"02", X"05", X"2c", X"23", X"aa", X"33", X"4c", X"3a", X"8d",
		X"52", X"0f", X"00", X"00", X"10", X"21", X"3c", X"05", X"00", X"3c", X"ae", X"c5", X"69", X"e2", X"f4",
		X"f2", X"00", X"00", X"52", X"41", X"1b", X"10", X"2d", X"a4", X"00", X"00", X"83", X"71", X"71", X"48",
		X"d7", X"bf", X"cd", X"ae", X"c7", X"d0", X"89", X"00", X"cf", X"af", X"ea", X"d2", X"f0", X"3a", X"23",
		X"1a", X"22", X"19", X"14", X"0c", X"38", X"3c", X"12", X"16", X"16", X"1a", X"2e", X"42", X"5e", X"4f",
		X"56", X"1e", X"10", X"12", X"1d", X"16", X"50", X"4d", X"39", X"1e", X"38", X"26", X"2d", X"46", X"4c",
		X"5b", X"02", X"04", X"09", X"12", X"01", X"03", X"04", X"00", X"00", X"7d", X"63", X"1a", X"02", X"00",
		X"00", X"07", X"06", X"06", X"1c", X"60", X"3e", X"04", X"16", X"1f", X"1d", X"f9", X"f9", X"d1", X"a4",
		X"ec", X"ef", X"a4", X"ce", X"ae", X"07", X"42", X"a8", X"00", X"07", X"8c", X"00", X"c1", X"ef", X"32",
		X"da", X"b9", X"97", X"cf", X"d8", X"ad", X"bd", X"4b", X"dc", X"cb", X"a8", X"e0", X"cd", X"80", X"00",
		X"27", X"14", X"03", X"2a", X"33", X"34", X"2c", X"17", X"0c", X"0a", X"0a", X"14", X"29", X"0a", X"21",
		X"22", X"3e", X"44", X"19", X"12", X"4e", X"56", X"55", X"45", X"51", X"31", X"25", X"23", X"53", X"5b",
		X"bf", X"d5", X"c2", X"9b", X"8f", X"63", X"93", X"bc", X"af", X"a1", X"c1", X"c2", X"a4", X"bf", X"ba",
		X"b1", X"c1", X"a5", X"b9", X"d3", X"bc", X"92", X"2f", X"12", X"1f", X"26", X"24", X"35", X"2b", X"21",
		X"2c", X"16", X"13", X"1a", X"11", X"18", X"08", X"6b", X"bb", X"d2", X"be", X"87", X"5e", X"61", X"4a",
		X"23", X"11", X"38", X"54", X"6a", X"62", X"4d", X"43", X"2e", X"28", X"20", X"38", X"42", X"40", X"2f",
		X"29", X"27", X"24", X"2e", X"2a", X"37", X"21", X"21", X"25", X"26", X"1e", X"24", X"27", X"2c", X"21",
		X"0d", X"0f", X"11", X"1a", X"24", X"24", X"1b", X"15", X"13", X"1c", X"15", X"1b", X"26", X"31", X"27",
		X"a7", X"bf", X"62", X"57", X"ac", X"88", X"96", X"d4", X"aa", X"56", X"8e", X"c4", X"d1", X"ac", X"8d",
		X"70", X"c8", X"97", X"88", X"cf", X"be", X"c6", X"ad", X"6a", X"32", X"19", X"0e", X"07", X"1c", X"28",
		X"23", X"27", X"21", X"18", X"1d", X"18", X"01", X"6a", X"c1", X"c7", X"c3", X"c6", X"bc", X"c3", X"bd",
		X"6a", X"38", X"5e", X"76", X"5a", X"49", X"3d", X"3f", X"46", X"34", X"2d", X"41", X"38", X"2d", X"2a",
		X"23", X"1d", X"26", X"33", X"36", X"3b", X"24", X"2f", X"32", X"2d", X"26", X"26", X"3a", X"3c", X"2f",
		X"16", X"1a", X"19", X"1e", X"1f", X"18", X"12", X"13", X"17", X"1b", X"13", X"25", X"41", X"27", X"28",
		X"8d", X"81", X"2f", X"af", X"ca", X"d9", X"c2", X"ab", X"88", X"35", X"35", X"88", X"77", X"b8", X"cd",
		X"54", X"9a", X"d6", X"c7", X"d0", X"b6", X"a2", X"be", X"aa", X"80", X"36", X"58", X"4b", X"1a", X"24",
		X"29", X"2a", X"2e", X"26", X"2f", X"21", X"0d", X"3f", X"83", X"a0", X"b4", X"c3", X"bc", X"b1", X"a3",
		X"7d", X"58", X"72", X"6a", X"5a", X"27", X"30", X"4e", X"48", X"2e", X"29", X"39", X"33", X"27", X"20",
		X"1f", X"1e", X"12", X"1b", X"1b", X"2a", X"2f", X"1a", X"30", X"26", X"21", X"2a", X"40", X"47", X"3e",
		X"1c", X"23", X"24", X"28", X"1c", X"15", X"12", X"16", X"1a", X"1f", X"19", X"2e", X"48", X"22", X"22",
		X"70", X"0c", X"3d", X"de", X"ce", X"c5", X"d2", X"bc", X"3e", X"00", X"0c", X"1b", X"08", X"73", X"91",
		X"31", X"17", X"bf", X"d4", X"c5", X"b9", X"b6", X"8d", X"6e", X"58", X"3a", X"8d", X"b2", X"86", X"3c",
		X"2e", X"2c", X"22", X"1e", X"27", X"20", X"1b", X"10", X"39", X"85", X"a2", X"a7", X"90", X"7e", X"72",
		X"3c", X"5e", X"69", X"6b", X"3b", X"20", X"2f", X"45", X"46", X"29", X"23", X"32", X"33", X"22", X"24",
		X"21", X"23", X"07", X"69", X"64", X"10", X"17", X"10", X"19", X"26", X"11", X"25", X"3f", X"48", X"44",
		X"1f", X"28", X"2b", X"30", X"20", X"0e", X"0f", X"17", X"18", X"1e", X"1f", X"2f", X"40", X"26", X"21",
		X"96", X"8c", X"7f", X"96", X"71", X"bb", X"db", X"a7", X"7a", X"65", X"22", X"08", X"14", X"95", X"66",
		X"63", X"51", X"24", X"65", X"dc", X"c2", X"d1", X"8f", X"95", X"94", X"82", X"4a", X"8f", X"ac", X"a4",
		X"7d", X"4c", X"19", X"18", X"2e", X"12", X"14", X"14", X"1b", X"6a", X"8e", X"aa", X"93", X"57", X"49",
		X"51", X"51", X"60", X"57", X"2c", X"37", X"49", X"48", X"35", X"27", X"27", X"3a", X"23", X"1b", X"50",
		X"5d", X"05", X"58", X"b1", X"bc", X"60", X"00", X"2c", X"19", X"1d", X"1c", X"22", X"42", X"4c", X"48",
		X"24", X"29", X"29", X"33", X"29", X"13", X"14", X"1a", X"19", X"1b", X"19", X"27", X"31", X"45", X"39",
		X"c7", X"ca", X"db", X"88", X"3a", X"7c", X"d3", X"ad", X"c5", X"bd", X"b0", X"6a", X"a4", X"b9", X"8a",
		X"8c", X"c4", X"c9", X"a5", X"d1", X"d8", X"a7", X"23", X"8d", X"ad", X"b2", X"7c", X"3f", X"60", X"6f",
		X"76", X"7e", X"3d", X"1b", X"28", X"13", X"19", X"1c", X"0e", X"7d", X"a1", X"c8", X"c2", X"61", X"4d",
		X"49", X"46", X"41", X"3f", X"34", X"3e", X"4a", X"47", X"30", X"32", X"32", X"24", X"26", X"1a", X"68",
		X"ac", X"74", X"7f", X"ad", X"bc", X"8d", X"20", X"3e", X"40", X"41", X"1c", X"18", X"3c", X"51", X"53",
		X"2a", X"24", X"2a", X"3a", X"34", X"27", X"19", X"16", X"17", X"18", X"11", X"19", X"1f", X"36", X"37",
		X"9d", X"90", X"b5", X"dc", X"8c", X"ab", X"c6", X"8b", X"c6", X"c7", X"93", X"aa", X"d1", X"bd", X"c1",
		X"8e", X"4a", X"8c", X"cb", X"92", X"b7", X"bf", X"73", X"45", X"96", X"af", X"8a", X"72", X"55", X"2d",
		X"67", X"70", X"5c", X"25", X"1a", X"2a", X"1f", X"1a", X"0d", X"62", X"af", X"c9", X"d8", X"7c", X"38",
		X"41", X"3e", X"44", X"42", X"33", X"4f", X"4b", X"47", X"51", X"38", X"23", X"2e", X"34", X"26", X"41",
		X"b5", X"c9", X"af", X"a8", X"b2", X"a5", X"83", X"8c", X"74", X"48", X"3a", X"39", X"3c", X"57", X"5d",
		X"3c", X"33", X"3b", X"47", X"41", X"31", X"1e", X"1a", X"1f", X"24", X"1d", X"1d", X"19", X"34", X"33",
		X"38", X"76", X"c6", X"cc", X"dd", X"d6", X"cb", X"bb", X"bd", X"d0", X"7b", X"91", X"dd", X"de", X"da",
		X"61", X"0b", X"c0", X"b3", X"ad", X"90", X"b5", X"e5", X"92", X"60", X"94", X"87", X"95", X"a5", X"8d",
		X"9b", X"c0", X"b5", X"40", X"32", X"a9", X"76", X"1c", X"05", X"33", X"cb", X"bb", X"c8", X"bd", X"82",
		X"3f", X"36", X"3c", X"27", X"4d", X"59", X"55", X"5f", X"61", X"3f", X"36", X"31", X"2c", X"32", X"1d",
		X"8f", X"c9", X"b5", X"d3", X"cc", X"cb", X"be", X"a2", X"7b", X"4a", X"38", X"49", X"4b", X"5d", X"62",
		X"52", X"50", X"54", X"54", X"4b", X"40", X"39", X"3d", X"3b", X"38", X"31", X"2b", X"1f", X"36", X"31",
		X"16", X"4f", X"c6", X"a7", X"a8", X"b6", X"c2", X"b7", X"ce", X"d3", X"5a", X"43", X"82", X"bc", X"d4",
		X"b4", X"90", X"ac", X"b1", X"d2", X"9e", X"50", X"76", X"7c", X"9b", X"98", X"b8", X"ad", X"be", X"b8",
		X"c5", X"cf", X"d5", X"41", X"39", X"a3", X"80", X"2e", X"60", X"57", X"c6", X"bb", X"ad", X"d4", X"c4",
		X"9e", X"6d", X"3c", X"32", X"4d", X"69", X"4e", X"45", X"43", X"47", X"4a", X"40", X"3c", X"2f", X"16",
		X"45", X"88", X"9b", X"c7", X"d6", X"d7", X"bd", X"a3", X"97", X"6e", X"42", X"45", X"4f", X"5e", X"62",
		X"67", X"6c", X"5a", X"5b", X"52", X"46", X"3c", X"3c", X"37", X"34", X"30", X"25", X"21", X"22", X"20",
		X"72", X"09", X"2b", X"3f", X"6a", X"93", X"a8", X"a6", X"b2", X"d0", X"44", X"70", X"6b", X"c5", X"a7",
		X"b4", X"ba", X"b4", X"8b", X"af", X"6a", X"cc", X"82", X"74", X"78", X"98", X"96", X"8d", X"a0", X"97",
		X"a7", X"b9", X"bf", X"41", X"32", X"74", X"27", X"32", X"80", X"71", X"86", X"be", X"c0", X"ba", X"c4",
		X"bd", X"c2", X"61", X"0f", X"30", X"64", X"82", X"63", X"22", X"54", X"4f", X"56", X"3c", X"21", X"15",
		X"19", X"4a", X"77", X"ab", X"c3", X"d2", X"bd", X"ad", X"96", X"78", X"39", X"33", X"3d", X"51", X"60",
		X"72", X"80", X"6e", X"63", X"52", X"3c", X"39", X"31", X"25", X"27", X"1e", X"16", X"20", X"1e", X"1c",
		X"60", X"41", X"34", X"28", X"35", X"59", X"63", X"99", X"ac", X"c7", X"48", X"88", X"cc", X"cc", X"cc",
		X"91", X"b5", X"b4", X"68", X"77", X"4d", X"3e", X"ad", X"6c", X"66", X"60", X"3f", X"3e", X"31", X"5c",
		X"ae", X"a0", X"9e", X"30", X"4c", X"ab", X"5b", X"69", X"70", X"a1", X"0c", X"4f", X"ba", X"b7", X"aa",
		X"ab", X"c5", X"ba", X"3c", X"7d", X"ac", X"c7", X"cb", X"4f", X"2d", X"4f", X"5b", X"4d", X"16", X"1a",
		X"1a", X"1a", X"46", X"90", X"bc", X"b6", X"7b", X"50", X"4a", X"37", X"32", X"22", X"1a", X"31", X"46",
		X"60", X"7c", X"7c", X"6f", X"54", X"34", X"1e", X"21", X"19", X"10", X"11", X"22", X"22", X"1b", X"1c",
		X"5e", X"3b", X"21", X"1b", X"46", X"48", X"6b", X"af", X"91", X"67", X"39", X"c5", X"a9", X"c9", X"c2",
		X"a7", X"6d", X"aa", X"b1", X"85", X"78", X"52", X"9b", X"71", X"54", X"3e", X"43", X"2a", X"08", X"4c",
		X"b4", X"b2", X"b5", X"1e", X"69", X"b8", X"a0", X"b6", X"bb", X"d2", X"6f", X"74", X"ae", X"ae", X"9a",
		X"ba", X"cc", X"d0", X"ca", X"a3", X"74", X"99", X"ab", X"89", X"32", X"48", X"48", X"4b", X"55", X"26",
		X"22", X"21", X"1c", X"22", X"51", X"52", X"3a", X"3e", X"51", X"5f", X"44", X"2b", X"03", X"14", X"28",
		X"48", X"6f", X"83", X"75", X"50", X"2d", X"21", X"22", X"1d", X"20", X"1c", X"24", X"27", X"1c", X"18",
		X"6d", X"3b", X"1e", X"0b", X"22", X"26", X"49", X"72", X"25", X"2e", X"4a", X"a6", X"6b", X"1d", X"92",
		X"92", X"88", X"91", X"da", X"a2", X"b5", X"c7", X"ad", X"7a", X"3f", X"50", X"2a", X"2a", X"20", X"59",
		X"a7", X"b4", X"a7", X"1f", X"67", X"d0", X"b2", X"c6", X"d1", X"ea", X"a4", X"72", X"84", X"9b", X"94",
		X"bc", X"be", X"b2", X"c6", X"c2", X"8c", X"ac", X"c0", X"9e", X"5c", X"47", X"54", X"60", X"52", X"4a",
		X"21", X"3e", X"3b", X"22", X"31", X"38", X"18", X"38", X"54", X"62", X"5d", X"33", X"0a", X"0c", X"17",
		X"37", X"5d", X"82", X"80", X"5e", X"2b", X"25", X"23", X"20", X"22", X"1f", X"28", X"2a", X"20", X"1b",
		X"75", X"39", X"0b", X"13", X"11", X"13", X"15", X"51", X"34", X"2b", X"4d", X"34", X"15", X"14", X"16",
		X"be", X"c7", X"a5", X"c5", X"ba", X"c9", X"c5", X"b1", X"64", X"37", X"1e", X"1d", X"6c", X"5b", X"3f",
		X"58", X"56", X"62", X"28", X"4f", X"bc", X"c4", X"b6", X"c1", X"b6", X"b1", X"54", X"57", X"7c", X"42",
		X"69", X"c3", X"a5", X"98", X"be", X"a2", X"a9", X"a3", X"7c", X"7a", X"5b", X"4d", X"4f", X"59", X"59",
		X"4c", X"55", X"61", X"3c", X"53", X"3f", X"26", X"1c", X"31", X"50", X"67", X"59", X"1e", X"21", X"33",
		X"46", X"54", X"7a", X"82", X"62", X"31", X"29", X"2b", X"2d", X"1d", X"1d", X"29", X"21", X"19", X"18",
		X"6a", X"44", X"1b", X"1e", X"23", X"1b", X"15", X"1d", X"22", X"1f", X"5f", X"25", X"33", X"1d", X"1d",
		X"90", X"e2", X"d1", X"cb", X"b7", X"44", X"a3", X"b9", X"bf", X"96", X"3b", X"3f", X"75", X"36", X"49",
		X"39", X"8e", X"ab", X"1a", X"4c", X"9c", X"a2", X"c9", X"94", X"8a", X"c3", X"95", X"7b", X"56", X"16",
		X"74", X"af", X"ae", X"aa", X"cb", X"8b", X"53", X"52", X"a7", X"9f", X"4d", X"4b", X"3a", X"2f", X"7b",
		X"80", X"59", X"80", X"7e", X"6a", X"4b", X"1a", X"25", X"1d", X"34", X"56", X"60", X"41", X"3d", X"4f",
		X"57", X"48", X"66", X"7b", X"69", X"3a", X"4b", X"43", X"48", X"46", X"3c", X"27", X"20", X"15", X"15",
		X"34", X"54", X"1b", X"20", X"1d", X"15", X"1c", X"21", X"1c", X"1a", X"58", X"26", X"1f", X"43", X"2a",
		X"13", X"76", X"a5", X"9f", X"b5", X"9d", X"a1", X"c5", X"b4", X"83", X"79", X"73", X"23", X"7d", X"ae",
		X"91", X"b5", X"bc", X"1a", X"78", X"c3", X"ba", X"bc", X"ae", X"9c", X"85", X"ac", X"b4", X"a9", X"26",
		X"74", X"a1", X"b6", X"bd", X"c1", X"ad", X"5d", X"61", X"a9", X"a7", X"54", X"28", X"36", X"15", X"6e",
		X"ab", X"7d", X"84", X"bb", X"a4", X"4f", X"18", X"21", X"1a", X"12", X"31", X"53", X"4e", X"4d", X"7c",
		X"a1", X"8b", X"92", X"95", X"81", X"4a", X"51", X"49", X"5a", X"57", X"5c", X"4a", X"36", X"15", X"12",
		X"16", X"5b", X"22", X"25", X"1b", X"1b", X"18", X"32", X"2a", X"23", X"60", X"21", X"0b", X"30", X"34",
		X"09", X"b4", X"e2", X"bc", X"d0", X"dd", X"95", X"98", X"54", X"3a", X"40", X"49", X"83", X"ab", X"ac",
		X"70", X"67", X"85", X"21", X"22", X"57", X"1c", X"64", X"d9", X"63", X"76", X"b6", X"b3", X"74", X"47",
		X"59", X"aa", X"ba", X"bf", X"94", X"ba", X"b7", X"89", X"50", X"82", X"4a", X"34", X"2d", X"21", X"41",
		X"96", X"9e", X"80", X"c3", X"b6", X"79", X"5d", X"58", X"0e", X"06", X"13", X"25", X"38", X"64", X"9f",
		X"b3", X"d4", X"cd", X"c5", X"d3", X"5f", X"27", X"49", X"3a", X"42", X"41", X"44", X"40", X"3c", X"33",
		X"36", X"2e", X"27", X"1b", X"39", X"50", X"34", X"1d", X"25", X"38", X"4c", X"6b", X"52", X"3c", X"2b",
		X"1c", X"6b", X"c0", X"67", X"63", X"6a", X"7c", X"8d", X"89", X"31", X"4c", X"22", X"48", X"7d", X"98",
		X"72", X"09", X"2c", X"4f", X"62", X"c6", X"ab", X"b4", X"d4", X"c5", X"bf", X"b2", X"c0", X"8f", X"68",
		X"24", X"57", X"d4", X"bd", X"c8", X"d2", X"ba", X"bf", X"8a", X"80", X"5c", X"56", X"41", X"24", X"1d",
		X"77", X"ba", X"b7", X"bc", X"b7", X"aa", X"8c", X"5a", X"15", X"03", X"00", X"07", X"1a", X"43", X"6b",
		X"8c", X"b3", X"c2", X"9b", X"c7", X"ae", X"26", X"14", X"2e", X"35", X"2e", X"2c", X"40", X"33", X"33",
		X"27", X"2b", X"21", X"14", X"26", X"50", X"29", X"49", X"20", X"49", X"45", X"6b", X"38", X"56", X"55",
		X"2b", X"38", X"5e", X"70", X"4e", X"45", X"c1", X"8e", X"b6", X"96", X"15", X"05", X"24", X"51", X"96",
		X"68", X"1c", X"36", X"5f", X"19", X"5b", X"fe", X"a7", X"f4", X"59", X"ec", X"ac", X"99", X"c0", X"e8",
		X"89", X"09", X"57", X"c8", X"ce", X"e5", X"b7", X"e2", X"f0", X"c6", X"78", X"57", X"2d", X"28", X"13",
		X"87", X"c8", X"ce", X"d3", X"af", X"90", X"3e", X"08", X"00", X"1c", X"66", X"6c", X"5c", X"7f", X"7c",
		X"85", X"6e", X"ad", X"a7", X"a3", X"d6", X"af", X"52", X"4e", X"45", X"35", X"18", X"28", X"33", X"34",
		X"14", X"23", X"24", X"21", X"03", X"60", X"21", X"9a", X"74", X"42", X"43", X"68", X"83", X"49", X"43",
		X"2f", X"29", X"36", X"3a", X"58", X"72", X"9f", X"f3", X"c2", X"b1", X"d0", X"32", X"00", X"31", X"21",
		X"0e", X"46", X"3c", X"3b", X"1f", X"01", X"30", X"c0", X"be", X"3c", X"ff", X"70", X"91", X"c1", X"7b",
		X"11", X"b6", X"a4", X"5e", X"b5", X"43", X"55", X"c8", X"c3", X"cd", X"c5", X"53", X"20", X"20", X"36",
		X"5b", X"ac", X"bf", X"b6", X"cb", X"9e", X"3d", X"00", X"04", X"44", X"a2", X"cb", X"b0", X"b1", X"b3",
		X"a9", X"6e", X"a6", X"de", X"c4", X"c1", X"bc", X"8e", X"5d", X"56", X"36", X"1a", X"17", X"35", X"37",
		X"3f", X"19", X"0c", X"0e", X"1f", X"60", X"38", X"a9", X"95", X"89", X"3d", X"2b", X"73", X"71", X"65",
		X"31", X"25", X"0a", X"44", X"ac", X"7c", X"1a", X"a3", X"cf", X"ea", X"b9", X"86", X"da", X"a0", X"c6",
		X"cd", X"2a", X"24", X"39", X"1a", X"20", X"1b", X"33", X"f3", X"38", X"c1", X"b7", X"98", X"45", X"0b",
		X"8f", X"bd", X"b8", X"c9", X"d4", X"d4", X"66", X"c2", X"c9", X"9f", X"43", X"6d", X"82", X"55", X"38",
		X"46", X"50", X"53", X"6f", X"97", X"a2", X"63", X"34", X"30", X"1e", X"59", X"bf", X"b6", X"b7", X"b2",
		X"ae", X"74", X"88", X"9f", X"be", X"cf", X"c1", X"9f", X"86", X"59", X"1f", X"18", X"17", X"3b", X"3e",
		X"26", X"32", X"12", X"48", X"b1", X"93", X"2f", X"a1", X"7d", X"bf", X"95", X"34", X"1b", X"39", X"4f",
		X"35", X"2c", X"55", X"95", X"a3", X"5a", X"56", X"a7", X"91", X"c5", X"e1", X"5a", X"b1", X"cc", X"c7",
		X"83", X"00", X"24", X"35", X"20", X"16", X"07", X"80", X"c5", X"4a", X"54", X"b5", X"6a", X"55", X"24",
		X"12", X"67", X"ba", X"d6", X"b0", X"e8", X"e0", X"bf", X"bd", X"ec", X"52", X"92", X"9c", X"84", X"5c",
		X"43", X"52", X"4f", X"67", X"77", X"7b", X"5e", X"4a", X"54", X"51", X"0b", X"4c", X"9e", X"c9", X"b9",
		X"69", X"7a", X"61", X"7c", X"7c", X"91", X"bd", X"89", X"8f", X"4a", X"1d", X"22", X"26", X"3f", X"40",
		X"26", X"20", X"16", X"21", X"ca", X"c2", X"37", X"b0", X"8a", X"bc", X"e2", X"d7", X"99", X"1d", X"72",
		X"2e", X"1a", X"a4", X"b6", X"ab", X"9c", X"86", X"d1", X"cf", X"bb", X"a2", X"4a", X"6e", X"cd", X"8e",
		X"03", X"0d", X"24", X"38", X"19", X"18", X"0c", X"26", X"ae", X"5a", X"14", X"db", X"81", X"72", X"1a",
		X"37", X"1e", X"02", X"37", X"00", X"c8", X"c5", X"c2", X"b1", X"bc", X"b0", X"45", X"62", X"a2", X"8b",
		X"73", X"2d", X"38", X"7f", X"95", X"99", X"87", X"4f", X"65", X"78", X"5d", X"41", X"af", X"c4", X"ac",
		X"a1", X"c3", X"5c", X"4b", X"4a", X"2f", X"3b", X"4b", X"48", X"2d", X"21", X"23", X"22", X"41", X"43",
		X"24", X"33", X"41", X"38", X"2c", X"8e", X"16", X"7d", X"5c", X"e6", X"ca", X"da", X"c6", X"55", X"28",
		X"36", X"23", X"a1", X"e3", X"a1", X"22", X"79", X"af", X"66", X"50", X"15", X"5a", X"2c", X"8f", X"de",
		X"7a", X"02", X"2b", X"34", X"24", X"09", X"3f", X"be", X"77", X"61", X"1b", X"9f", X"a3", X"e9", X"7b",
		X"17", X"20", X"10", X"38", X"40", X"2f", X"3f", X"65", X"b1", X"a8", X"b7", X"34", X"8f", X"de", X"bd",
		X"72", X"4d", X"91", X"93", X"95", X"a9", X"81", X"84", X"56", X"8a", X"7d", X"6b", X"ae", X"ab", X"8a",
		X"a2", X"bc", X"64", X"2b", X"37", X"32", X"1c", X"34", X"2a", X"29", X"24", X"22", X"22", X"43", X"42",
		X"16", X"31", X"69", X"8d", X"3e", X"80", X"d5", X"bc", X"9c", X"7a", X"e8", X"cd", X"c3", X"94", X"2e",
		X"35", X"20", X"6b", X"d1", X"9e", X"1e", X"b7", X"e8", X"91", X"00", X"6a", X"73", X"65", X"18", X"9a",
		X"90", X"a8", X"46", X"2c", X"00", X"3a", X"b4", X"c1", X"8a", X"55", X"32", X"7d", X"90", X"ce", X"c4",
		X"73", X"aa", X"88", X"05", X"c0", X"25", X"41", X"4b", X"45", X"a5", X"9b", X"c8", X"7e", X"c4", X"e8",
		X"98", X"b1", X"8c", X"59", X"88", X"6d", X"65", X"69", X"62", X"9a", X"8e", X"55", X"52", X"61", X"66",
		X"6a", X"87", X"85", X"25", X"2d", X"2d", X"25", X"20", X"2a", X"1e", X"21", X"24", X"18", X"19", X"25",
		X"19", X"10", X"0b", X"1d", X"79", X"a3", X"a1", X"b7", X"c7", X"cc", X"36", X"77", X"ff", X"77", X"d0",
		X"38", X"29", X"4f", X"b4", X"69", X"2d", X"bc", X"d3", X"95", X"04", X"96", X"ab", X"7d", X"ab", X"a6",
		X"90", X"82", X"7b", X"3b", X"cc", X"6e", X"43", X"9b", X"eb", X"58", X"36", X"8a", X"65", X"b8", X"de",
		X"97", X"98", X"9b", X"73", X"c6", X"b1", X"9c", X"93", X"6b", X"40", X"34", X"ba", X"99", X"d9", X"b3",
		X"fe", X"6c", X"4b", X"7e", X"8d", X"3c", X"65", X"3b", X"6c", X"7a", X"7e", X"4a", X"33", X"26", X"3d",
		X"34", X"92", X"8c", X"39", X"22", X"23", X"26", X"1b", X"1a", X"21", X"22", X"1a", X"1d", X"29", X"25",
		X"3b", X"0f", X"1b", X"23", X"1c", X"81", X"aa", X"ba", X"d7", X"e8", X"b8", X"6a", X"19", X"73", X"c3",
		X"40", X"34", X"2d", X"66", X"1a", X"22", X"68", X"a3", X"30", X"4f", X"cd", X"9c", X"c7", X"aa", X"a2",
		X"c3", X"c0", X"4c", X"8b", X"d7", X"ad", X"7e", X"97", X"33", X"66", X"23", X"8b", X"ed", X"b4", X"c4",
		X"a9", X"5e", X"21", X"69", X"58", X"79", X"93", X"65", X"3d", X"2a", X"26", X"10", X"32", X"eb", X"d0",
		X"6d", X"5d", X"73", X"b4", X"1f", X"4d", X"5a", X"59", X"49", X"40", X"31", X"40", X"2f", X"46", X"54",
		X"45", X"4d", X"71", X"2d", X"28", X"20", X"21", X"1c", X"1b", X"32", X"2d", X"18", X"1f", X"27", X"28",
		X"9f", X"36", X"00", X"19", X"00", X"00", X"5b", X"af", X"b6", X"cd", X"af", X"5b", X"00", X"a6", X"ee",
		X"41", X"28", X"19", X"10", X"63", X"02", X"23", X"40", X"04", X"4c", X"38", X"f4", X"91", X"d1", X"be",
		X"bf", X"e9", X"df", X"b5", X"d3", X"e0", X"78", X"0a", X"4f", X"6d", X"3b", X"5f", X"e6", X"c3", X"92",
		X"b4", X"4d", X"20", X"20", X"6e", X"a7", X"5b", X"38", X"2d", X"27", X"18", X"33", X"29", X"5d", X"73",
		X"77", X"4a", X"db", X"a9", X"60", X"5c", X"57", X"40", X"20", X"26", X"17", X"1a", X"20", X"4d", X"67",
		X"62", X"38", X"3c", X"30", X"32", X"30", X"21", X"24", X"25", X"3e", X"36", X"1d", X"21", X"27", X"2a",
		X"c1", X"75", X"00", X"04", X"09", X"1a", X"00", X"84", X"d7", X"99", X"d2", X"00", X"3a", X"e1", X"53",
		X"47", X"2d", X"23", X"0b", X"2b", X"3e", X"0c", X"69", X"1f", X"2e", X"0c", X"5e", X"eb", X"ac", X"b1",
		X"c3", X"db", X"e3", X"b5", X"b4", X"e0", X"9a", X"4d", X"32", X"6e", X"35", X"38", X"c5", X"c1", X"6e",
		X"56", X"1c", X"44", X"2e", X"bc", X"ae", X"85", X"20", X"2e", X"22", X"29", X"2d", X"1f", X"49", X"6d",
		X"61", X"8e", X"db", X"ce", X"88", X"72", X"4f", X"29", X"56", X"42", X"25", X"30", X"2b", X"4c", X"5d",
		X"56", X"67", X"38", X"59", X"35", X"37", X"22", X"23", X"26", X"41", X"3d", X"2a", X"3c", X"15", X"21",
		X"98", X"53", X"0d", X"0b", X"02", X"24", X"00", X"99", X"c6", X"de", X"43", X"06", X"96", X"b4", X"8b",
		X"36", X"3a", X"25", X"0d", X"1c", X"46", X"3c", X"14", X"0e", X"4f", X"9a", X"5b", X"83", X"ad", X"89",
		X"a8", X"6f", X"d7", X"b9", X"a1", X"cf", X"d7", X"9d", X"59", X"47", X"53", X"40", X"64", X"9a", X"61",
		X"01", X"6f", X"75", X"1a", X"4e", X"a4", X"5b", X"11", X"14", X"49", X"56", X"48", X"00", X"55", X"82",
		X"66", X"a6", X"fe", X"c3", X"7c", X"9b", X"2e", X"32", X"5a", X"4b", X"32", X"1e", X"23", X"4b", X"59",
		X"65", X"51", X"64", X"42", X"56", X"32", X"28", X"24", X"27", X"45", X"42", X"2e", X"4c", X"24", X"20",
		X"64", X"27", X"0e", X"10", X"0c", X"1a", X"2d", X"e2", X"c5", X"fe", X"09", X"21", X"e3", X"a7", X"85",
		X"74", X"2d", X"2f", X"0d", X"28", X"49", X"29", X"2a", X"2b", X"76", X"8e", X"a9", X"da", X"a1", X"d7",
		X"fe", X"e6", X"d6", X"c5", X"ee", X"ee", X"d8", X"a5", X"64", X"47", X"4c", X"35", X"89", X"a9", X"0a",
		X"8d", X"52", X"7a", X"43", X"08", X"81", X"61", X"22", X"4a", X"7a", X"63", X"37", X"29", X"96", X"6b",
		X"69", X"2c", X"c1", X"be", X"bc", X"bd", X"3d", X"14", X"2b", X"35", X"4d", X"38", X"0a", X"6d", X"aa",
		X"88", X"71", X"54", X"55", X"33", X"28", X"24", X"24", X"2f", X"4a", X"4c", X"35", X"44", X"22", X"25",
		X"89", X"68", X"12", X"0a", X"1c", X"19", X"18", X"00", X"20", X"0e", X"1d", X"57", X"90", X"71", X"63",
		X"29", X"49", X"22", X"29", X"21", X"3c", X"3b", X"11", X"1c", X"4c", X"83", X"4a", X"54", X"5d", X"48",
		X"2c", X"a3", X"be", X"48", X"58", X"ed", X"b1", X"a7", X"7b", X"55", X"67", X"11", X"a4", X"e4", X"a6",
		X"80", X"40", X"81", X"36", X"0b", X"49", X"5e", X"62", X"52", X"4e", X"66", X"02", X"aa", X"6d", X"71",
		X"2b", X"2e", X"06", X"ba", X"d3", X"b6", X"44", X"24", X"18", X"25", X"38", X"35", X"1e", X"44", X"bf",
		X"cb", X"b3", X"59", X"43", X"33", X"2b", X"20", X"22", X"34", X"44", X"51", X"3b", X"2f", X"25", X"27",
		X"61", X"2b", X"47", X"0e", X"1d", X"13", X"23", X"2d", X"1f", X"22", X"09", X"a1", X"d9", X"4b", X"55",
		X"0f", X"5b", X"1a", X"32", X"28", X"3b", X"53", X"1a", X"30", X"19", X"1c", X"22", X"06", X"3f", X"46",
		X"15", X"93", X"c9", X"86", X"6d", X"c2", X"e3", X"bd", X"a0", X"7c", X"81", X"3c", X"a9", X"d4", X"d8",
		X"d2", X"a8", X"ab", X"8c", X"bd", X"00", X"99", X"81", X"2a", X"3f", X"17", X"4b", X"b4", X"5e", X"4c",
		X"22", X"65", X"6f", X"41", X"a2", X"b7", X"94", X"6a", X"20", X"15", X"2e", X"26", X"23", X"20", X"71",
		X"b2", X"d9", X"99", X"4c", X"2e", X"21", X"23", X"2a", X"36", X"46", X"50", X"34", X"16", X"17", X"2c",
		X"56", X"4e", X"1a", X"39", X"08", X"1a", X"65", X"1e", X"18", X"2f", X"0f", X"a6", X"3c", X"69", X"66",
		X"0d", X"57", X"1f", X"3a", X"22", X"21", X"67", X"03", X"a3", X"7d", X"23", X"2b", X"12", X"4a", X"33",
		X"1b", X"f8", X"be", X"7d", X"c5", X"ee", X"d9", X"d2", X"a0", X"63", X"89", X"ff", X"b1", X"7f", X"ff",
		X"dc", X"de", X"b9", X"5e", X"6b", X"71", X"47", X"75", X"95", X"13", X"0b", X"9c", X"80", X"2d", X"1b",
		X"1e", X"37", X"a8", X"85", X"9c", X"a6", X"ab", X"b3", X"58", X"00", X"19", X"11", X"88", X"87", X"b8",
		X"a2", X"c0", X"b8", X"9b", X"27", X"15", X"21", X"26", X"39", X"49", X"49", X"3e", X"2d", X"2b", X"29",
		X"3f", X"7e", X"15", X"2e", X"12", X"2d", X"54", X"1f", X"30", X"1a", X"2a", X"15", X"09", X"45", X"2a",
		X"43", X"4a", X"2d", X"38", X"2b", X"16", X"2b", X"2f", X"87", X"9c", X"1a", X"25", X"1a", X"35", X"5e",
		X"5b", X"4b", X"9b", X"aa", X"b2", X"cb", X"9e", X"d2", X"b7", X"66", X"03", X"e2", X"ed", X"ff", X"3b",
		X"0c", X"c6", X"ea", X"37", X"4f", X"26", X"a7", X"a0", X"e3", X"07", X"30", X"00", X"0a", X"10", X"53",
		X"38", X"50", X"4d", X"c4", X"c9", X"96", X"3e", X"5a", X"51", X"0e", X"27", X"3e", X"28", X"6e", X"39",
		X"4e", X"bb", X"cc", X"c5", X"a8", X"39", X"0f", X"1f", X"35", X"44", X"4f", X"5a", X"76", X"24", X"2a",
		X"47", X"7f", X"74", X"0d", X"1e", X"5c", X"9b", X"1c", X"16", X"3b", X"23", X"18", X"3c", X"42", X"07",
		X"00", X"7d", X"4f", X"21", X"28", X"2a", X"3f", X"20", X"19", X"0b", X"3b", X"3f", X"4f", X"47", X"13",
		X"88", X"af", X"bc", X"3e", X"ff", X"ed", X"85", X"0a", X"05", X"0d", X"43", X"3b", X"63", X"5a", X"ff",
		X"ad", X"dc", X"46", X"71", X"41", X"e0", X"43", X"92", X"3c", X"5d", X"3c", X"26", X"14", X"36", X"53",
		X"8e", X"80", X"83", X"95", X"8b", X"b8", X"be", X"56", X"62", X"5a", X"08", X"15", X"44", X"8b", X"85",
		X"d0", X"aa", X"b6", X"c7", X"a7", X"8b", X"24", X"2d", X"2d", X"27", X"58", X"82", X"8b", X"2b", X"24",
		X"69", X"55", X"59", X"91", X"14", X"20", X"50", X"46", X"16", X"85", X"7d", X"38", X"3a", X"1b", X"22",
		X"ba", X"dc", X"84", X"22", X"29", X"20", X"0e", X"71", X"73", X"28", X"36", X"53", X"1a", X"32", X"08",
		X"45", X"73", X"84", X"3a", X"4a", X"fa", X"8c", X"0a", X"32", X"1a", X"13", X"5a", X"2a", X"42", X"f0",
		X"e7", X"5d", X"cf", X"ef", X"90", X"9b", X"3e", X"19", X"8b", X"84", X"7f", X"5e", X"3b", X"40", X"53",
		X"61", X"4b", X"1f", X"9b", X"9f", X"a8", X"db", X"6f", X"17", X"28", X"2f", X"24", X"2e", X"2f", X"12",
		X"29", X"28", X"7b", X"a0", X"b0", X"7b", X"37", X"2e", X"1f", X"17", X"2c", X"60", X"6e", X"53", X"6c",
		X"65", X"5f", X"07", X"5d", X"80", X"11", X"2a", X"07", X"84", X"88", X"82", X"51", X"30", X"50", X"93",
		X"84", X"bc", X"4f", X"21", X"2e", X"3c", X"42", X"6b", X"b6", X"7a", X"24", X"92", X"21", X"0a", X"40",
		X"2d", X"33", X"1b", X"66", X"0a", X"1f", X"8b", X"10", X"22", X"38", X"0b", X"30", X"3a", X"7d", X"ff",
		X"21", X"77", X"da", X"bc", X"dc", X"6a", X"0c", X"41", X"64", X"49", X"7a", X"49", X"61", X"2c", X"28",
		X"28", X"0a", X"2c", X"6c", X"5c", X"81", X"e0", X"00", X"a4", X"60", X"13", X"1f", X"29", X"25", X"26",
		X"28", X"24", X"42", X"6b", X"b0", X"82", X"20", X"17", X"1a", X"14", X"23", X"55", X"4a", X"6c", X"65",
		X"61", X"20", X"24", X"03", X"6f", X"78", X"12", X"20", X"98", X"e5", X"a5", X"bc", X"9f", X"78", X"69",
		X"5a", X"aa", X"50", X"21", X"1d", X"43", X"3f", X"41", X"4b", X"42", X"33", X"21", X"38", X"14", X"55",
		X"00", X"14", X"23", X"7d", X"55", X"30", X"01", X"16", X"28", X"39", X"18", X"38", X"39", X"08", X"2a",
		X"a1", X"48", X"00", X"0f", X"95", X"18", X"46", X"67", X"43", X"5c", X"45", X"4a", X"aa", X"1c", X"1c",
		X"0b", X"0b", X"2c", X"33", X"0a", X"64", X"9d", X"3a", X"c6", X"ae", X"57", X"1a", X"21", X"2b", X"1c",
		X"1f", X"1a", X"19", X"37", X"7d", X"7d", X"34", X"30", X"28", X"27", X"25", X"4c", X"4f", X"65", X"66",
		X"97", X"1e", X"1c", X"2d", X"1c", X"95", X"2f", X"23", X"23", X"ff", X"cd", X"be", X"ae", X"f2", X"62",
		X"76", X"94", X"60", X"3b", X"16", X"31", X"17", X"5f", X"0e", X"17", X"19", X"08", X"19", X"33", X"00",
		X"1a", X"00", X"69", X"92", X"66", X"00", X"0e", X"58", X"2a", X"66", X"40", X"10", X"16", X"31", X"34",
		X"35", X"15", X"33", X"8f", X"13", X"3d", X"58", X"64", X"42", X"3d", X"5a", X"59", X"02", X"2a", X"1a",
		X"16", X"1b", X"28", X"2f", X"31", X"3c", X"2c", X"58", X"79", X"8d", X"77", X"34", X"1b", X"24", X"11",
		X"04", X"13", X"18", X"07", X"21", X"42", X"2d", X"35", X"54", X"56", X"13", X"31", X"46", X"62", X"68",
		X"b4", X"ff", X"4f", X"22", X"32", X"00", X"13", X"39", X"79", X"3b", X"da", X"cb", X"a5", X"7b", X"fb",
		X"ad", X"df", X"86", X"90", X"76", X"3f", X"16", X"54", X"11", X"40", X"d0", X"b3", X"46", X"03", X"17",
		X"33", X"b3", X"a4", X"72", X"00", X"91", X"d0", X"be", X"a9", X"28", X"2c", X"24", X"2c", X"25", X"52",
		X"3c", X"06", X"0e", X"52", X"b2", X"1d", X"6c", X"25", X"1e", X"70", X"5c", X"3a", X"12", X"40", X"3f",
		X"40", X"4f", X"53", X"4c", X"4d", X"48", X"42", X"21", X"41", X"5d", X"99", X"47", X"5d", X"46", X"3b",
		X"32", X"29", X"2c", X"5a", X"2e", X"29", X"21", X"2d", X"4c", X"4d", X"27", X"39", X"3f", X"1c", X"0d",
		X"53", X"98", X"cc", X"0a", X"69", X"79", X"1d", X"13", X"90", X"d0", X"d5", X"e8", X"47", X"57", X"68",
		X"dd", X"c0", X"75", X"48", X"5b", X"64", X"1d", X"37", X"55", X"0d", X"7b", X"e9", X"c4", X"9b", X"0b",
		X"9d", X"82", X"9d", X"a0", X"00", X"d6", X"e5", X"b0", X"c1", X"69", X"2a", X"33", X"26", X"51", X"63",
		X"7e", X"70", X"3a", X"09", X"5d", X"00", X"5d", X"1d", X"5c", X"66", X"44", X"3c", X"14", X"3c", X"32",
		X"45", X"4f", X"2f", X"34", X"20", X"19", X"40", X"61", X"08", X"2e", X"49", X"73", X"c4", X"82", X"61",
		X"55", X"58", X"7d", X"62", X"5a", X"40", X"2d", X"39", X"5d", X"4b", X"2e", X"2c", X"4a", X"0e", X"06",
		X"60", X"53", X"90", X"0e", X"92", X"cf", X"db", X"8d", X"a5", X"bc", X"c6", X"e9", X"55", X"75", X"c5",
		X"c1", X"de", X"95", X"77", X"36", X"39", X"33", X"21", X"4d", X"23", X"0a", X"97", X"e9", X"c4", X"ba",
		X"a9", X"47", X"e5", X"3b", X"37", X"b3", X"a3", X"df", X"db", X"b3", X"18", X"34", X"32", X"46", X"40",
		X"5a", X"6c", X"3e", X"21", X"21", X"1b", X"3a", X"13", X"52", X"b6", X"b5", X"ac", X"1c", X"28", X"1f",
		X"20", X"1d", X"7c", X"4e", X"29", X"32", X"22", X"14", X"0b", X"50", X"a1", X"9a", X"b8", X"bc", X"83",
		X"5f", X"7f", X"52", X"77", X"45", X"3b", X"12", X"47", X"7b", X"57", X"2c", X"2c", X"42", X"06", X"0b",
		X"13", X"2b", X"1b", X"20", X"1d", X"80", X"ca", X"df", X"db", X"9f", X"8c", X"d5", X"ec", X"ea", X"a8",
		X"d4", X"92", X"53", X"34", X"34", X"17", X"25", X"1a", X"2e", X"3a", X"ca", X"d1", X"c0", X"e3", X"bf",
		X"e1", X"ff", X"1d", X"1b", X"09", X"35", X"b8", X"ad", X"a4", X"03", X"34", X"0a", X"3e", X"3e", X"4f",
		X"6f", X"27", X"2f", X"10", X"13", X"55", X"31", X"21", X"74", X"ff", X"c7", X"58", X"6b", X"c1", X"db",
		X"6a", X"63", X"c0", X"90", X"65", X"1d", X"15", X"14", X"31", X"2b", X"65", X"d5", X"bc", X"cf", X"d1",
		X"64", X"63", X"70", X"53", X"3b", X"24", X"05", X"2c", X"75", X"44", X"2a", X"30", X"3a", X"0f", X"06",
		X"2a", X"72", X"28", X"41", X"10", X"00", X"9c", X"c1", X"ee", X"d3", X"d9", X"d3", X"f2", X"c0", X"8a",
		X"c6", X"a6", X"18", X"40", X"30", X"07", X"37", X"27", X"0c", X"73", X"a0", X"b5", X"c3", X"ba", X"65",
		X"a0", X"cf", X"00", X"0f", X"00", X"6d", X"80", X"a4", X"ae", X"07", X"21", X"9a", X"60", X"53", X"89",
		X"1e", X"13", X"71", X"17", X"1f", X"56", X"50", X"b0", X"f6", X"43", X"0c", X"00", X"49", X"b1", X"92",
		X"f6", X"59", X"df", X"d5", X"8a", X"0f", X"37", X"65", X"34", X"4a", X"53", X"38", X"f3", X"d4", X"d5",
		X"69", X"76", X"99", X"99", X"89", X"8c", X"77", X"7d", X"45", X"4a", X"0a", X"44", X"1d", X"22", X"0d",
		X"67", X"57", X"41", X"4a", X"4d", X"85", X"6f", X"da", X"c3", X"92", X"b9", X"d7", X"d7", X"64", X"94",
		X"7f", X"db", X"0d", X"3f", X"26", X"10", X"10", X"3a", X"14", X"22", X"4d", X"8f", X"da", X"d0", X"ac",
		X"a6", X"d7", X"cf", X"1f", X"00", X"78", X"66", X"7c", X"a7", X"3e", X"98", X"5f", X"67", X"92", X"9a",
		X"0a", X"8c", X"9c", X"85", X"4b", X"b8", X"ba", X"75", X"05", X"14", X"56", X"cb", X"08", X"d6", X"a0",
		X"96", X"cb", X"a2", X"e8", X"af", X"0c", X"38", X"34", X"48", X"9d", X"96", X"b6", X"c3", X"e4", X"76",
		X"4a", X"bd", X"ca", X"99", X"51", X"3a", X"3e", X"49", X"4a", X"48", X"0d", X"47", X"34", X"0e", X"0f",
		X"29", X"2f", X"56", X"8a", X"c5", X"bc", X"af", X"91", X"d8", X"69", X"9c", X"90", X"c3", X"b2", X"5c",
		X"62", X"9c", X"11", X"37", X"22", X"14", X"0a", X"08", X"1e", X"29", X"29", X"29", X"60", X"7b", X"93",
		X"d2", X"bd", X"e1", X"dc", X"00", X"32", X"cb", X"b5", X"c1", X"df", X"59", X"62", X"86", X"39", X"ae",
		X"be", X"a2", X"a9", X"3e", X"2c", X"5a", X"31", X"18", X"17", X"57", X"f6", X"56", X"a5", X"c0", X"ea",
		X"d8", X"bf", X"c1", X"e8", X"58", X"20", X"3b", X"44", X"85", X"b8", X"aa", X"b7", X"e9", X"fa", X"72",
		X"0d", X"b2", X"c3", X"ad", X"a5", X"6c", X"25", X"04", X"57", X"47", X"1c", X"33", X"48", X"0d", X"07",
		X"65", X"30", X"8c", X"60", X"b1", X"d1", X"c2", X"c3", X"fb", X"2b", X"5e", X"e1", X"a3", X"d7", X"b7",
		X"1f", X"13", X"23", X"1b", X"20", X"12", X"10", X"3c", X"13", X"30", X"2a", X"7d", X"5a", X"94", X"6f",
		X"c6", X"ba", X"a2", X"af", X"45", X"00", X"f9", X"c9", X"d6", X"ef", X"a8", X"91", X"8f", X"4b", X"1e",
		X"db", X"d0", X"bd", X"0c", X"40", X"31", X"6b", X"64", X"3b", X"3a", X"e3", X"7c", X"31", X"84", X"7e",
		X"ae", X"d6", X"00", X"74", X"71", X"0e", X"74", X"8a", X"58", X"5e", X"74", X"7d", X"58", X"72", X"ff",
		X"84", X"d0", X"d7", X"a0", X"00", X"09", X"00", X"1c", X"52", X"48", X"16", X"28", X"3e", X"09", X"08",
		X"6a", X"5b", X"84", X"5f", X"47", X"dd", X"da", X"bb", X"c9", X"e6", X"eb", X"b1", X"de", X"c0", X"85",
		X"14", X"15", X"18", X"1f", X"0c", X"17", X"00", X"5b", X"21", X"2b", X"3a", X"bf", X"5e", X"a5", X"3a",
		X"ac", X"aa", X"89", X"00", X"84", X"ab", X"be", X"c7", X"46", X"8e", X"fc", X"c2", X"83", X"b4", X"ee",
		X"9c", X"d7", X"cf", X"03", X"57", X"70", X"54", X"12", X"9f", X"db", X"a2", X"9a", X"63", X"50", X"bc",
		X"22", X"c8", X"00", X"cb", X"c8", X"6a", X"52", X"8d", X"61", X"3f", X"3f", X"68", X"0e", X"14", X"dd",
		X"bd", X"de", X"9c", X"ec", X"24", X"00", X"02", X"19", X"5b", X"55", X"17", X"1d", X"2b", X"30", X"7c",
		X"45", X"8d", X"75", X"63", X"5a", X"ba", X"13", X"98", X"df", X"c9", X"ae", X"bc", X"a3", X"d2", X"00",
		X"14", X"20", X"12", X"21", X"27", X"25", X"16", X"0c", X"25", X"22", X"98", X"b1", X"c9", X"77", X"2e",
		X"86", X"80", X"97", X"b5", X"b5", X"c2", X"e8", X"a8", X"48", X"06", X"ac", X"c2", X"6c", X"7d", X"8e",
		X"b3", X"ac", X"e1", X"82", X"29", X"39", X"03", X"9f", X"8c", X"bb", X"c9", X"6e", X"af", X"57", X"3e",
		X"37", X"cf", X"e8", X"a8", X"a0", X"6e", X"32", X"37", X"5a", X"6a", X"8c", X"41", X"13", X"64", X"ce",
		X"cc", X"b8", X"5e", X"ad", X"fe", X"3a", X"27", X"19", X"51", X"38", X"23", X"21", X"2c", X"7a", X"78",
		X"74", X"74", X"60", X"5d", X"16", X"4f", X"47", X"97", X"ca", X"e7", X"c7", X"dc", X"87", X"d1", X"3a",
		X"00", X"14", X"2b", X"39", X"38", X"32", X"1c", X"29", X"26", X"1f", X"31", X"4f", X"11", X"3f", X"51",
		X"5f", X"90", X"3a", X"8e", X"a4", X"c0", X"af", X"d3", X"5f", X"c8", X"cf", X"cb", X"87", X"82", X"a0",
		X"6b", X"2a", X"c6", X"f3", X"45", X"06", X"2f", X"50", X"7d", X"f3", X"a2", X"3e", X"05", X"1f", X"04",
		X"47", X"ae", X"9e", X"b9", X"a1", X"65", X"6d", X"74", X"74", X"89", X"58", X"15", X"64", X"12", X"89",
		X"f4", X"46", X"1f", X"4c", X"d4", X"79", X"79", X"59", X"36", X"26", X"2c", X"31", X"1e", X"78", X"7b",
		X"38", X"25", X"2d", X"61", X"43", X"22", X"14", X"19", X"d7", X"c5", X"4b", X"5a", X"c5", X"8d", X"71",
		X"1d", X"2b", X"1e", X"10", X"24", X"09", X"21", X"10", X"1a", X"25", X"14", X"15", X"32", X"42", X"29",
		X"09", X"1d", X"6c", X"6d", X"b6", X"a6", X"9f", X"96", X"ec", X"aa", X"ab", X"8e", X"73", X"67", X"1b",
		X"2b", X"24", X"23", X"d4", X"78", X"08", X"39", X"4a", X"24", X"fa", X"08", X"05", X"11", X"0b", X"1b",
		X"2d", X"96", X"9b", X"d9", X"50", X"63", X"6d", X"8a", X"ab", X"54", X"07", X"42", X"1b", X"31", X"46",
		X"71", X"27", X"27", X"27", X"74", X"dd", X"43", X"46", X"37", X"49", X"40", X"38", X"3c", X"78", X"77",
		X"3f", X"1d", X"11", X"5f", X"6f", X"00", X"1a", X"0f", X"1e", X"a8", X"2e", X"61", X"32", X"bc", X"79",
		X"5c", X"0b", X"14", X"1a", X"18", X"15", X"0d", X"13", X"07", X"36", X"1a", X"20", X"30", X"33", X"30",
		X"18", X"39", X"03", X"12", X"ff", X"ec", X"b6", X"cb", X"92", X"e9", X"ab", X"95", X"56", X"0b", X"02",
		X"e7", X"c8", X"00", X"b4", X"00", X"29", X"3f", X"3b", X"1b", X"07", X"22", X"29", X"03", X"12", X"3b",
		X"23", X"74", X"80", X"bf", X"2d", X"50", X"69", X"ac", X"92", X"20", X"87", X"4b", X"30", X"35", X"4a",
		X"23", X"22", X"41", X"3d", X"1b", X"5f", X"12", X"3e", X"44", X"41", X"35", X"3a", X"3e", X"68", X"99",
		X"42", X"04", X"09", X"04", X"5d", X"3a", X"05", X"0e", X"49", X"74", X"52", X"20", X"c9", X"88", X"8b",
		X"67", X"05", X"13", X"39", X"0d", X"13", X"16", X"0b", X"10", X"2f", X"13", X"0f", X"3d", X"56", X"05",
		X"10", X"44", X"0d", X"3a", X"f1", X"de", X"fd", X"b7", X"68", X"fa", X"ce", X"c3", X"80", X"0e", X"a0",
		X"9a", X"af", X"0f", X"47", X"22", X"25", X"51", X"1d", X"37", X"16", X"34", X"08", X"0c", X"17", X"09",
		X"1e", X"43", X"4f", X"5b", X"2d", X"3f", X"92", X"88", X"08", X"73", X"7a", X"21", X"39", X"2c", X"2d",
		X"2c", X"0c", X"18", X"27", X"76", X"05", X"96", X"3d", X"34", X"2a", X"2c", X"22", X"37", X"95", X"98",
		X"10", X"1c", X"0d", X"03", X"04", X"2a", X"06", X"1a", X"42", X"5c", X"69", X"89", X"dd", X"c2", X"63",
		X"7b", X"5a", X"05", X"1f", X"15", X"03", X"0a", X"18", X"0c", X"15", X"16", X"21", X"46", X"00", X"02",
		X"2c", X"09", X"11", X"11", X"55", X"b3", X"52", X"0c", X"14", X"5d", X"bc", X"b9", X"53", X"1a", X"ae",
		X"82", X"d5", X"ed", X"56", X"ba", X"84", X"56", X"6f", X"e1", X"66", X"07", X"0b", X"0e", X"0f", X"3a",
		X"59", X"1b", X"3f", X"9b", X"2b", X"63", X"62", X"11", X"6a", X"4e", X"30", X"3e", X"31", X"1d", X"17",
		X"38", X"da", X"af", X"b8", X"2f", X"5e", X"20", X"29", X"2c", X"2a", X"37", X"2e", X"22", X"98", X"96",
		X"19", X"0d", X"15", X"10", X"0f", X"06", X"0a", X"1b", X"4f", X"52", X"53", X"21", X"62", X"9b", X"73",
		X"6a", X"20", X"1c", X"1a", X"11", X"24", X"04", X"11", X"0b", X"0f", X"7e", X"e2", X"6f", X"bc", X"17",
		X"1d", X"35", X"28", X"1d", X"1d", X"58", X"1e", X"d6", X"38", X"01", X"00", X"91", X"b6", X"a9", X"aa",
		X"aa", X"ad", X"4e", X"50", X"40", X"d4", X"7b", X"3d", X"93", X"dd", X"15", X"09", X"00", X"54", X"7b",
		X"28", X"31", X"57", X"3b", X"3e", X"41", X"1f", X"3a", X"6d", X"57", X"20", X"1b", X"1b", X"23", X"27",
		X"7a", X"51", X"30", X"0f", X"33", X"22", X"27", X"34", X"29", X"2e", X"27", X"2c", X"33", X"90", X"96",
		X"22", X"20", X"0a", X"03", X"0b", X"0b", X"01", X"2e", X"51", X"48", X"69", X"3e", X"46", X"05", X"24",
		X"84", X"77", X"07", X"20", X"09", X"09", X"05", X"16", X"06", X"29", X"c9", X"38", X"dd", X"fd", X"de",
		X"03", X"0e", X"12", X"13", X"57", X"2e", X"16", X"b2", X"f7", X"27", X"0a", X"55", X"d3", X"95", X"b1",
		X"ce", X"a2", X"9e", X"8b", X"ce", X"d1", X"45", X"23", X"c5", X"a1", X"b8", X"d4", X"b0", X"06", X"2f",
		X"1f", X"21", X"33", X"18", X"29", X"1b", X"3e", X"4b", X"3f", X"3b", X"57", X"51", X"50", X"3c", X"3d",
		X"27", X"28", X"22", X"23", X"1e", X"16", X"1a", X"21", X"16", X"30", X"27", X"19", X"22", X"33", X"44",
		X"0a", X"0a", X"14", X"06", X"06", X"09", X"03", X"0a", X"3b", X"34", X"b8", X"36", X"47", X"3b", X"8e",
		X"57", X"19", X"09", X"0c", X"1d", X"2b", X"3d", X"0d", X"01", X"46", X"b9", X"d1", X"76", X"ec", X"f5",
		X"fa", X"01", X"02", X"53", X"3c", X"1c", X"11", X"31", X"a8", X"00", X"06", X"84", X"6c", X"72", X"49",
		X"db", X"c3", X"cb", X"b2", X"cc", X"d5", X"8c", X"00", X"d3", X"af", X"e8", X"d6", X"f5", X"3f", X"26",
		X"19", X"26", X"19", X"12", X"14", X"44", X"44", X"1d", X"21", X"1e", X"22", X"36", X"4a", X"6a", X"57",
		X"61", X"29", X"18", X"1a", X"25", X"11", X"56", X"5a", X"41", X"1e", X"31", X"1e", X"28", X"46", X"48",
		X"62", X"0d", X"13", X"12", X"12", X"08", X"09", X"07", X"03", X"08", X"8c", X"6c", X"1a", X"09", X"03",
		X"00", X"0d", X"11", X"11", X"25", X"66", X"41", X"0a", X"1f", X"25", X"28", X"ff", X"ff", X"d7", X"a7",
		X"f2", X"f8", X"b2", X"d1", X"ad", X"09", X"47", X"b1", X"00", X"08", X"9a", X"03", X"c0", X"f1", X"37",
		X"e3", X"bf", X"98", X"d8", X"e3", X"b9", X"c7", X"53", X"e7", X"cf", X"a9", X"e9", X"d8", X"8c", X"06",
		X"2f", X"1f", X"07", X"2b", X"3e", X"40", X"37", X"23", X"1a", X"18", X"18", X"22", X"34", X"16", X"2c",
		X"2e", X"4c", X"52", X"27", X"20", X"52", X"66", X"6b", X"56", X"5b", X"32", X"24", X"25", X"48", X"49",
		X"ec", X"de", X"b4", X"96", X"a9", X"95", X"bb", X"d4", X"dc", X"aa", X"b3", X"bd", X"be", X"f1", X"e2",
		X"c9", X"c1", X"bd", X"d8", X"e7", X"9e", X"93", X"0c", X"00", X"1f", X"3e", X"43", X"49", X"0d", X"22",
		X"09", X"00", X"00", X"03", X"18", X"30", X"1c", X"93", X"d3", X"9f", X"a9", X"70", X"65", X"79", X"5e",
		X"4b", X"29", X"05", X"20", X"3f", X"3d", X"25", X"1f", X"13", X"19", X"19", X"04", X"17", X"1b", X"07",
		X"05", X"0c", X"15", X"27", X"2e", X"32", X"1b", X"0a", X"00", X"15", X"14", X"00", X"2b", X"27", X"1b",
		X"00", X"00", X"00", X"10", X"00", X"09", X"03", X"00", X"01", X"0d", X"09", X"0f", X"1c", X"16", X"0f",
		X"b9", X"cc", X"6b", X"68", X"b9", X"8e", X"af", X"fe", X"bc", X"63", X"97", X"d5", X"de", X"b2", X"a6",
		X"9a", X"da", X"bc", X"b3", X"f4", X"dd", X"f5", X"bc", X"61", X"44", X"3e", X"39", X"2c", X"3b", X"57",
		X"32", X"1e", X"0c", X"00", X"17", X"30", X"2e", X"99", X"cb", X"99", X"ae", X"ac", X"b6", X"db", X"ea",
		X"99", X"42", X"30", X"3d", X"42", X"31", X"0f", X"15", X"33", X"27", X"1c", X"08", X"20", X"15", X"00",
		X"00", X"0a", X"19", X"22", X"2a", X"34", X"1f", X"0e", X"00", X"02", X"14", X"0e", X"2e", X"35", X"2a",
		X"00", X"00", X"00", X"0c", X"07", X"05", X"02", X"05", X"0b", X"12", X"0d", X"1f", X"3e", X"11", X"16",
		X"a8", X"7a", X"0f", X"c9", X"f7", X"db", X"d4", X"d7", X"a3", X"2e", X"15", X"a2", X"a4", X"ba", X"df",
		X"80", X"b6", X"f8", X"e7", X"f0", X"de", X"c7", X"ec", X"cd", X"9c", X"58", X"78", X"6b", X"42", X"49",
		X"57", X"4d", X"20", X"15", X"20", X"2e", X"38", X"55", X"62", X"58", X"a6", X"b2", X"ad", X"be", X"ce",
		X"93", X"37", X"2a", X"3d", X"34", X"06", X"0c", X"2a", X"3b", X"3c", X"41", X"0c", X"0d", X"06", X"00",
		X"00", X"11", X"20", X"33", X"2e", X"26", X"1d", X"00", X"00", X"00", X"00", X"0f", X"53", X"43", X"2c",
		X"00", X"00", X"00", X"00", X"01", X"00", X"00", X"06", X"0d", X"12", X"0e", X"22", X"3f", X"13", X"16",
		X"72", X"1f", X"39", X"f9", X"ed", X"bd", X"e7", X"e0", X"40", X"12", X"08", X"36", X"27", X"6b", X"a6",
		X"55", X"36", X"d9", X"d9", X"e4", X"db", X"cd", X"bb", X"a4", X"77", X"54", X"92", X"d1", X"a8", X"53",
		X"5c", X"62", X"1c", X"1d", X"2a", X"2c", X"37", X"1c", X"1c", X"4c", X"9c", X"a6", X"93", X"8a", X"8e",
		X"48", X"41", X"30", X"43", X"05", X"00", X"08", X"14", X"32", X"45", X"4b", X"0a", X"00", X"00", X"00",
		X"00", X"0f", X"23", X"91", X"8e", X"27", X"13", X"00", X"00", X"00", X"00", X"00", X"69", X"5f", X"40",
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"05", X"06", X"16", X"26", X"1a", X"17",
		X"92", X"ae", X"94", X"c2", X"89", X"98", X"dc", X"d3", X"76", X"87", X"37", X"34", X"2c", X"72", X"67",
		X"8f", X"77", X"4c", X"68", X"ff", X"f2", X"ff", X"bf", X"b6", X"ba", X"aa", X"4d", X"be", X"dc", X"df",
		X"ad", X"6d", X"15", X"28", X"4d", X"2b", X"2a", X"36", X"3c", X"75", X"8a", X"ba", X"b2", X"70", X"5f",
		X"73", X"72", X"6b", X"1f", X"0d", X"1d", X"1d", X"1a", X"24", X"2c", X"2a", X"02", X"04", X"01", X"24",
		X"2f", X"00", X"5d", X"b4", X"c9", X"7c", X"0c", X"0b", X"00", X"00", X"00", X"00", X"4f", X"68", X"56",
		X"03", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"09", X"13", X"32", X"29",
		X"a2", X"e2", X"e7", X"89", X"43", X"81", X"eb", X"cc", X"a0", X"d5", X"bc", X"6b", X"ad", X"be", X"a2",
		X"ab", X"e3", X"ff", X"bb", X"f9", X"ea", X"e0", X"4b", X"a9", X"cc", X"e8", X"92", X"67", X"72", X"a8",
		X"9e", X"9a", X"39", X"35", X"54", X"2c", X"25", X"3e", X"40", X"a4", X"9d", X"e2", X"ee", X"7a", X"59",
		X"6b", X"78", X"68", X"64", X"6d", X"49", X"1d", X"1b", X"0c", X"1a", X"41", X"49", X"5f", X"25", X"3b",
		X"80", X"50", X"67", X"bc", X"c1", X"7f", X"00", X"17", X"1a", X"05", X"00", X"00", X"41", X"43", X"31",
		X"03", X"00", X"00", X"00", X"00", X"07", X"00", X"00", X"00", X"00", X"00", X"00", X"04", X"28", X"2b",
		X"65", X"88", X"ab", X"ce", X"8a", X"a2", X"c8", X"b3", X"8e", X"bf", X"89", X"9c", X"cf", X"b4", X"c3",
		X"b6", X"60", X"ab", X"e6", X"aa", X"b2", X"cd", X"80", X"6b", X"ac", X"ce", X"a5", X"8a", X"50", X"3b",
		X"74", X"96", X"55", X"3d", X"39", X"39", X"31", X"32", X"29", X"86", X"a8", X"e1", X"f7", X"8b", X"4a",
		X"59", X"5a", X"68", X"4e", X"50", X"65", X"55", X"52", X"55", X"42", X"4d", X"3a", X"51", X"3c", X"4b",
		X"c0", X"cd", X"b9", X"d2", X"cc", X"8a", X"3b", X"5b", X"61", X"1e", X"00", X"0f", X"56", X"3c", X"15",
		X"0b", X"20", X"11", X"07", X"17", X"10", X"00", X"00", X"04", X"0a", X"03", X"03", X"00", X"2b", X"2d",
		X"0f", X"77", X"c5", X"af", X"c2", X"b6", X"a9", X"bf", X"94", X"d1", X"7a", X"74", X"c2", X"be", X"b8",
		X"65", X"2a", X"bb", X"c3", X"d0", X"b1", X"ba", X"da", X"b0", X"7f", X"8f", X"97", X"b8", X"c6", X"92",
		X"90", X"de", X"a4", X"52", X"41", X"bb", X"a6", X"44", X"1f", X"6a", X"ba", X"cd", X"d7", X"cf", X"b2",
		X"67", X"50", X"73", X"4f", X"6d", X"7b", X"57", X"34", X"51", X"55", X"40", X"59", X"4c", X"54", X"1f",
		X"64", X"b9", X"cb", X"dd", X"e8", X"d3", X"97", X"65", X"57", X"2f", X"12", X"23", X"67", X"65", X"3b",
		X"15", X"2c", X"39", X"2e", X"25", X"16", X"12", X"1a", X"19", X"17", X"0f", X"09", X"00", X"30", X"2e",
		X"43", X"58", X"b8", X"a2", X"c2", X"e8", X"ea", X"cf", X"fb", X"dc", X"4c", X"3e", X"9c", X"ee", X"fc",
		X"cc", X"90", X"c4", X"d0", X"e6", X"80", X"51", X"53", X"63", X"9b", X"b0", X"d7", X"c1", X"a0", X"b9",
		X"a2", X"b6", X"c0", X"2a", X"40", X"bb", X"94", X"56", X"78", X"24", X"b1", X"a4", X"b4", X"ec", X"d8",
		X"c6", X"85", X"09", X"00", X"22", X"44", X"26", X"21", X"28", X"38", X"43", X"0c", X"11", X"0a", X"00",
		X"21", X"6d", X"8c", X"c0", X"da", X"d2", X"b7", X"8c", X"71", X"5d", X"38", X"1d", X"53", X"59", X"5c",
		X"50", X"46", X"49", X"51", X"2a", X"2b", X"24", X"26", X"25", X"25", X"24", X"19", X"17", X"07", X"08",
		X"84", X"16", X"34", X"50", X"77", X"99", X"c1", X"d0", X"c4", X"dd", X"4d", X"81", X"78", X"cb", X"c0",
		X"de", X"cc", X"d9", X"b6", X"d4", X"89", X"fb", X"91", X"6b", X"8a", X"bd", X"c1", X"b2", X"bf", X"c6",
		X"b6", X"b0", X"aa", X"27", X"2c", X"8c", X"54", X"61", X"8a", X"43", X"71", X"a4", X"ba", X"d2", X"f1",
		X"ec", X"cc", X"33", X"00", X"18", X"4c", X"54", X"39", X"0f", X"47", X"3e", X"1d", X"24", X"09", X"00",
		X"00", X"37", X"6a", X"9a", X"b7", X"cb", X"b8", X"8c", X"58", X"4d", X"27", X"1b", X"31", X"4a", X"5b",
		X"51", X"42", X"43", X"51", X"3a", X"29", X"29", X"23", X"19", X"1e", X"18", X"10", X"1d", X"08", X"0a",
		X"7b", X"3a", X"14", X"42", X"62", X"5b", X"75", X"c5", X"c7", X"c0", X"28", X"a2", X"f9", X"ce", X"de",
		X"bd", X"d1", X"d6", X"88", X"97", X"75", X"63", X"db", X"8f", X"82", X"82", X"5f", X"5e", X"59", X"81",
		X"dc", X"c3", X"90", X"1f", X"3d", X"b8", X"86", X"7f", X"4f", X"59", X"00", X"3e", X"ab", X"c4", X"d5",
		X"c1", X"a4", X"72", X"0f", X"57", X"8b", X"a3", X"a7", X"42", X"3b", X"67", X"2e", X"27", X"00", X"00",
		X"00", X"0d", X"54", X"a8", X"cf", X"b2", X"69", X"2d", X"0f", X"00", X"0a", X"07", X"2d", X"2d", X"34",
		X"3d", X"41", X"41", X"47", X"39", X"1f", X"0b", X"11", X"0c", X"03", X"06", X"16", X"19", X"0c", X"10",
		X"60", X"4e", X"1d", X"36", X"65", X"40", X"80", X"d3", X"93", X"7a", X"35", X"e0", X"c8", X"c1", X"d7",
		X"cb", X"8c", X"c4", X"b6", X"a4", X"9a", X"69", X"c9", X"a7", X"73", X"58", X"48", X"49", X"2a", X"63",
		X"e2", X"e8", X"af", X"1d", X"6c", X"c4", X"bc", X"c2", X"9e", X"99", X"69", X"73", X"b1", X"ba", X"b6",
		X"c6", X"af", X"97", X"a2", X"6d", X"48", X"72", X"7a", X"75", X"4e", X"70", X"20", X"15", X"29", X"00",
		X"00", X"0d", X"38", X"4a", X"7b", X"69", X"36", X"1f", X"1d", X"25", X"0f", X"00", X"2d", X"2b", X"24",
		X"29", X"3b", X"49", X"40", X"1b", X"0b", X"01", X"04", X"02", X"07", X"03", X"0b", X"0d", X"10", X"0e",
		X"69", X"5d", X"33", X"37", X"3a", X"03", X"4a", X"9e", X"21", X"50", X"5f", X"d2", X"83", X"00", X"93",
		X"be", X"ae", X"b9", X"dd", X"d1", X"e5", X"ff", X"dd", X"9b", X"65", X"78", X"2d", X"59", X"50", X"94",
		X"d7", X"d5", X"a3", X"2f", X"86", X"e9", X"c8", X"e8", X"f2", X"f5", X"a0", X"82", X"a3", X"b4", X"aa",
		X"de", X"df", X"bd", X"8e", X"a3", X"72", X"80", X"92", X"8d", X"61", X"4a", X"1c", X"41", X"38", X"1e",
		X"00", X"2d", X"40", X"25", X"3e", X"54", X"26", X"17", X"18", X"27", X"21", X"00", X"17", X"28", X"25",
		X"16", X"21", X"47", X"44", X"1b", X"05", X"00", X"01", X"01", X"04", X"01", X"0a", X"0c", X"0d", X"0b",
		X"50", X"51", X"17", X"14", X"1a", X"18", X"2d", X"70", X"0f", X"43", X"59", X"35", X"1e", X"19", X"2e",
		X"dd", X"e6", X"db", X"db", X"e2", X"db", X"fe", X"d9", X"80", X"56", X"54", X"33", X"94", X"6d", X"78",
		X"80", X"72", X"5e", X"42", X"7b", X"d5", X"d0", X"d8", X"f3", X"dd", X"ad", X"6e", X"83", X"95", X"4e",
		X"8b", X"f5", X"cc", X"bd", X"f7", X"ad", X"7c", X"77", X"58", X"62", X"6a", X"72", X"88", X"64", X"2c",
		X"20", X"31", X"49", X"4b", X"58", X"31", X"04", X"00", X"0b", X"14", X"20", X"21", X"23", X"13", X"11",
		X"1f", X"2e", X"3e", X"3b", X"2a", X"11", X"0a", X"0e", X"13", X"05", X"05", X"0e", X"06", X"0b", X"0c",
		X"32", X"3c", X"11", X"10", X"21", X"12", X"17", X"45", X"00", X"17", X"55", X"17", X"31", X"14", X"1f",
		X"b8", X"f8", X"f0", X"e6", X"cf", X"3f", X"b1", X"c6", X"e5", X"ac", X"5a", X"5a", X"8d", X"31", X"57",
		X"46", X"b4", X"a4", X"32", X"6b", X"ab", X"b4", X"e1", X"b0", X"ae", X"bc", X"ad", X"9a", X"65", X"28",
		X"8c", X"cb", X"d2", X"b6", X"e8", X"a1", X"5d", X"5d", X"ab", X"a9", X"77", X"57", X"57", X"45", X"85",
		X"8b", X"5d", X"8a", X"a8", X"84", X"30", X"00", X"00", X"0a", X"0a", X"16", X"36", X"5b", X"22", X"07",
		X"26", X"35", X"3c", X"3b", X"3f", X"19", X"2b", X"27", X"2d", X"2c", X"22", X"0d", X"05", X"0c", X"0f",
		X"0b", X"55", X"1a", X"03", X"02", X"00", X"00", X"25", X"00", X"1b", X"57", X"09", X"04", X"23", X"08",
		X"17", X"95", X"a0", X"af", X"d8", X"be", X"a6", X"ba", X"d2", X"a2", X"74", X"83", X"46", X"9e", X"b3",
		X"86", X"d3", X"ab", X"2c", X"87", X"d5", X"ea", X"e4", X"c8", X"d3", X"74", X"be", X"c3", X"bb", X"56",
		X"9c", X"bb", X"ed", X"e5", X"e1", X"cf", X"5f", X"36", X"99", X"bd", X"5e", X"50", X"56", X"37", X"70",
		X"80", X"6d", X"9a", X"c5", X"c0", X"57", X"00", X"00", X"00", X"00", X"0b", X"2d", X"6a", X"55", X"55",
		X"64", X"67", X"77", X"6f", X"5b", X"20", X"2a", X"26", X"38", X"36", X"3a", X"28", X"14", X"0f", X"0f",
		X"00", X"37", X"28", X"08", X"0d", X"0d", X"23", X"15", X"0b", X"00", X"66", X"04", X"00", X"22", X"3f",
		X"00", X"c8", X"f8", X"d0", X"e7", X"b7", X"88", X"ab", X"54", X"4e", X"56", X"5d", X"9a", X"85", X"9f",
		X"83", X"67", X"5f", X"37", X"37", X"89", X"47", X"81", X"ff", X"a2", X"50", X"cc", X"c8", X"a6", X"72",
		X"76", X"d1", X"f9", X"ea", X"be", X"d6", X"c3", X"87", X"37", X"92", X"5c", X"5f", X"57", X"3d", X"4d",
		X"94", X"85", X"90", X"d5", X"d8", X"9d", X"5d", X"50", X"00", X"18", X"18", X"21", X"5a", X"88", X"9f",
		X"ab", X"c5", X"df", X"ca", X"cf", X"44", X"06", X"22", X"11", X"19", X"18", X"17", X"0e", X"21", X"12",
		X"25", X"09", X"44", X"35", X"41", X"48", X"5f", X"29", X"14", X"13", X"69", X"85", X"5a", X"34", X"56",
		X"28", X"5b", X"da", X"89", X"8d", X"88", X"7c", X"73", X"7e", X"21", X"66", X"44", X"72", X"9b", X"98",
		X"58", X"00", X"0f", X"58", X"62", X"c0", X"ae", X"d7", X"ec", X"de", X"a2", X"bb", X"c0", X"89", X"6b",
		X"47", X"6f", X"ed", X"d9", X"c1", X"ee", X"d9", X"d0", X"64", X"8c", X"76", X"72", X"3a", X"40", X"3c",
		X"88", X"94", X"c3", X"d6", X"be", X"b6", X"97", X"65", X"18", X"12", X"09", X"01", X"21", X"4f", X"76",
		X"97", X"b6", X"d1", X"a5", X"c1", X"b2", X"1d", X"00", X"0b", X"0d", X"02", X"00", X"10", X"0c", X"0a",
		X"13", X"12", X"2e", X"20", X"38", X"4a", X"37", X"3c", X"0c", X"30", X"52", X"77", X"4a", X"50", X"63",
		X"1e", X"2b", X"4f", X"7f", X"7b", X"58", X"bd", X"ba", X"dc", X"89", X"06", X"14", X"51", X"64", X"92",
		X"94", X"42", X"10", X"51", X"24", X"60", X"f9", X"be", X"f3", X"72", X"c6", X"9e", X"a4", X"c5", X"e3",
		X"a0", X"08", X"70", X"f0", X"dd", X"f6", X"df", X"f5", X"fc", X"b9", X"6d", X"7f", X"3c", X"39", X"3b",
		X"9a", X"d4", X"c1", X"c8", X"c5", X"82", X"3f", X"1c", X"13", X"28", X"7e", X"81", X"72", X"71", X"7d",
		X"99", X"82", X"b9", X"bf", X"b8", X"f5", X"bd", X"48", X"2f", X"1d", X"06", X"00", X"00", X"0a", X"0b",
		X"00", X"1c", X"34", X"2c", X"26", X"7d", X"44", X"97", X"53", X"3b", X"53", X"73", X"a6", X"66", X"66",
		X"2c", X"2d", X"49", X"46", X"6e", X"7b", X"77", X"ff", X"c5", X"b5", X"e3", X"3e", X"14", X"3a", X"00",
		X"21", X"49", X"10", X"20", X"1b", X"00", X"22", X"cb", X"b0", X"44", X"da", X"55", X"8d", X"bc", X"6d",
		X"1c", X"a8", X"ac", X"6a", X"cc", X"5b", X"86", X"c6", X"ef", X"cc", X"cb", X"5f", X"37", X"38", X"67",
		X"59", X"d8", X"be", X"bc", X"f8", X"97", X"47", X"12", X"19", X"47", X"b6", X"c5", X"dd", X"aa", X"bd",
		X"bb", X"83", X"a9", X"f2", X"be", X"b6", X"aa", X"74", X"3e", X"3c", X"23", X"0b", X"0b", X"08", X"05",
		X"36", X"2e", X"3e", X"40", X"37", X"6c", X"5e", X"a0", X"8c", X"9e", X"6f", X"5d", X"8b", X"7d", X"8b",
		X"28", X"1c", X"1f", X"4a", X"9e", X"90", X"1e", X"c7", X"ff", X"e1", X"ce", X"8c", X"cc", X"b4", X"ca",
		X"f1", X"5c", X"1a", X"5d", X"45", X"26", X"00", X"38", X"ff", X"51", X"b7", X"db", X"c3", X"4b", X"00",
		X"94", X"d0", X"d1", X"da", X"d6", X"e2", X"7c", X"ba", X"dc", X"9e", X"4a", X"7e", X"84", X"63", X"4e",
		X"3e", X"63", X"52", X"76", X"91", X"8b", X"6f", X"3a", X"32", X"1b", X"65", X"9b", X"b0", X"a0", X"be",
		X"b4", X"76", X"85", X"ab", X"9a", X"b4", X"a5", X"81", X"6b", X"41", X"0a", X"00", X"00", X"3f", X"35",
		X"04", X"2b", X"15", X"66", X"c9", X"97", X"45", X"a3", X"5b", X"b8", X"98", X"52", X"33", X"3d", X"65",
		X"37", X"11", X"3a", X"a0", X"a6", X"72", X"88", X"d3", X"b4", X"aa", X"c6", X"65", X"b4", X"e4", X"f9",
		X"af", X"20", X"45", X"5b", X"34", X"0f", X"00", X"91", X"cf", X"38", X"75", X"db", X"7e", X"4e", X"08",
		X"23", X"71", X"a8", X"d6", X"c9", X"d5", X"c6", X"ab", X"c0", X"c1", X"47", X"92", X"b5", X"71", X"42",
		X"2f", X"55", X"24", X"5c", X"68", X"56", X"4d", X"42", X"3c", X"28", X"00", X"31", X"8f", X"a4", X"a8",
		X"61", X"62", X"38", X"63", X"61", X"5e", X"8d", X"5e", X"6f", X"31", X"06", X"07", X"06", X"26", X"1d",
		X"04", X"25", X"05", X"2b", X"e9", X"cb", X"40", X"ae", X"68", X"c1", X"d1", X"e1", X"b8", X"26", X"7b",
		X"2c", X"00", X"80", X"88", X"8c", X"a1", X"a8", X"e6", X"e8", X"96", X"7e", X"1c", X"4f", X"d2", X"b0",
		X"18", X"26", X"39", X"47", X"3b", X"24", X"00", X"3c", X"b6", X"64", X"29", X"ea", X"a3", X"7e", X"03",
		X"4d", X"26", X"0c", X"08", X"12", X"aa", X"b2", X"9e", X"9b", X"8e", X"c6", X"16", X"77", X"84", X"78",
		X"4f", X"17", X"0a", X"95", X"b8", X"95", X"66", X"37", X"40", X"4c", X"2b", X"17", X"d2", X"c0", X"8b",
		X"89", X"9e", X"30", X"19", X"20", X"0e", X"18", X"25", X"20", X"07", X"00", X"00", X"00", X"19", X"17",
		X"00", X"29", X"36", X"42", X"2e", X"92", X"3b", X"84", X"1b", X"dc", X"bf", X"e4", X"c8", X"59", X"4d",
		X"3d", X"00", X"97", X"a5", X"ae", X"58", X"a1", X"d0", X"74", X"2c", X"0b", X"1c", X"39", X"c5", X"ff",
		X"9b", X"10", X"1f", X"28", X"3e", X"00", X"00", X"dd", X"90", X"84", X"0f", X"93", X"bd", X"c9", X"3c",
		X"36", X"39", X"33", X"43", X"28", X"14", X"50", X"55", X"78", X"90", X"ba", X"3f", X"77", X"c3", X"ce",
		X"62", X"14", X"79", X"96", X"a2", X"b2", X"58", X"58", X"44", X"b1", X"7f", X"39", X"bb", X"b4", X"61",
		X"76", X"aa", X"8b", X"2d", X"05", X"13", X"00", X"04", X"00", X"00", X"00", X"00", X"00", X"15", X"12",
		X"00", X"0d", X"6f", X"70", X"30", X"72", X"e0", X"9f", X"7d", X"56", X"ee", X"b0", X"b5", X"86", X"39",
		X"18", X"34", X"81", X"e5", X"b5", X"00", X"aa", X"fb", X"91", X"12", X"80", X"87", X"7c", X"00", X"8d",
		X"a3", X"a8", X"20", X"42", X"12", X"6c", X"df", X"de", X"b1", X"94", X"0c", X"93", X"a5", X"ff", X"ef",
		X"90", X"d1", X"c7", X"30", X"ea", X"41", X"4d", X"49", X"2c", X"b5", X"ad", X"f3", X"a8", X"e0", X"f4",
		X"96", X"98", X"9c", X"6b", X"aa", X"91", X"65", X"61", X"53", X"ac", X"93", X"51", X"74", X"85", X"66",
		X"62", X"78", X"97", X"2a", X"29", X"12", X"04", X"00", X"01", X"00", X"00", X"00", X"00", X"00", X"04",
		X"08", X"00", X"28", X"37", X"81", X"9b", X"cc", X"c3", X"b6", X"a7", X"53", X"91", X"ff", X"6f", X"fb",
		X"44", X"19", X"69", X"d6", X"93", X"4b", X"bc", X"b9", X"8a", X"00", X"b0", X"cd", X"a7", X"c9", X"a6",
		X"76", X"77", X"5e", X"44", X"cc", X"68", X"46", X"be", X"ff", X"71", X"19", X"93", X"65", X"b2", X"e1",
		X"ba", X"b0", X"b4", X"8f", X"bf", X"cd", X"bb", X"a4", X"45", X"4c", X"4e", X"d6", X"92", X"f5", X"d2",
		X"ff", X"46", X"57", X"98", X"94", X"48", X"70", X"46", X"6f", X"89", X"88", X"44", X"3a", X"32", X"48",
		X"3f", X"95", X"9b", X"43", X"1c", X"27", X"1d", X"02", X"00", X"00", X"00", X"00", X"00", X"02", X"00",
		X"27", X"00", X"28", X"2f", X"2e", X"7b", X"b8", X"ad", X"c3", X"cf", X"c5", X"76", X"2b", X"6d", X"d1",
		X"33", X"27", X"1e", X"75", X"47", X"35", X"64", X"cf", X"56", X"42", X"be", X"ab", X"f4", X"bd", X"9e",
		X"ef", X"e6", X"26", X"7d", X"e2", X"b2", X"79", X"ae", X"32", X"7f", X"00", X"7d", X"f8", X"b9", X"bf",
		X"c0", X"5d", X"3a", X"91", X"67", X"8a", X"bb", X"78", X"49", X"1d", X"1b", X"38", X"41", X"fc", X"f8",
		X"80", X"69", X"66", X"a9", X"35", X"3f", X"5b", X"6d", X"5d", X"4c", X"49", X"55", X"45", X"38", X"55",
		X"59", X"61", X"7d", X"45", X"3d", X"3f", X"2f", X"12", X"00", X"0a", X"00", X"00", X"00", X"00", X"00",
		X"7e", X"2f", X"10", X"24", X"21", X"19", X"7e", X"ac", X"95", X"c6", X"bf", X"66", X"1e", X"c3", X"ff",
		X"3e", X"2c", X"2c", X"1c", X"79", X"0b", X"00", X"53", X"07", X"50", X"4b", X"ff", X"a7", X"da", X"96",
		X"d2", X"ec", X"b3", X"9a", X"cf", X"db", X"6a", X"15", X"41", X"75", X"0f", X"44", X"e2", X"be", X"84",
		X"bf", X"3f", X"28", X"2c", X"85", X"bf", X"8c", X"36", X"59", X"26", X"1e", X"3f", X"40", X"75", X"a4",
		X"75", X"76", X"da", X"af", X"8d", X"55", X"61", X"52", X"35", X"29", X"2b", X"14", X"4d", X"46", X"71",
		X"74", X"4d", X"3f", X"44", X"2c", X"25", X"0f", X"0a", X"06", X"24", X"23", X"0e", X"15", X"00", X"00",
		X"b8", X"8a", X"30", X"36", X"21", X"26", X"22", X"7b", X"ce", X"ae", X"ff", X"2b", X"52", X"ed", X"79",
		X"3e", X"24", X"38", X"11", X"1d", X"52", X"10", X"8d", X"51", X"25", X"21", X"64", X"dd", X"c0", X"b5",
		X"e7", X"ff", X"d9", X"d9", X"df", X"e6", X"77", X"52", X"45", X"87", X"2b", X"5c", X"f0", X"c7", X"4b",
		X"5b", X"2f", X"5d", X"3f", X"be", X"bc", X"9b", X"18", X"41", X"21", X"30", X"3e", X"21", X"57", X"83",
		X"59", X"a1", X"da", X"d5", X"82", X"5b", X"5b", X"2f", X"58", X"3f", X"31", X"0c", X"25", X"35", X"69",
		X"5c", X"69", X"35", X"65", X"11", X"1c", X"06", X"05", X"0b", X"29", X"28", X"11", X"1e", X"19", X"18",
		X"76", X"4c", X"10", X"29", X"1a", X"28", X"14", X"9b", X"a4", X"d7", X"46", X"24", X"ae", X"b8", X"a1",
		X"38", X"1f", X"0a", X"18", X"1f", X"5e", X"6e", X"40", X"31", X"34", X"7f", X"66", X"86", X"c5", X"bb",
		X"d4", X"92", X"f8", X"df", X"b5", X"c8", X"bb", X"ae", X"63", X"35", X"74", X"66", X"78", X"93", X"45",
		X"12", X"79", X"63", X"1a", X"67", X"91", X"41", X"00", X"17", X"1e", X"4b", X"48", X"17", X"42", X"68",
		X"52", X"a9", X"d3", X"b8", X"6d", X"76", X"1d", X"2a", X"42", X"22", X"19", X"03", X"14", X"26", X"48",
		X"5d", X"39", X"3b", X"29", X"3b", X"00", X"00", X"00", X"07", X"2c", X"2b", X"13", X"2c", X"0b", X"00",
		X"42", X"2c", X"00", X"1a", X"2b", X"23", X"36", X"e0", X"a3", X"ff", X"00", X"2b", X"ff", X"b0", X"8e",
		X"72", X"08", X"0b", X"00", X"09", X"4e", X"4b", X"3f", X"44", X"51", X"6a", X"7b", X"bb", X"a6", X"f9",
		X"ff", X"ff", X"eb", X"d4", X"ff", X"fa", X"c1", X"bb", X"6c", X"51", X"61", X"44", X"ab", X"b5", X"00",
		X"a3", X"5a", X"84", X"14", X"1d", X"63", X"4e", X"00", X"34", X"4c", X"79", X"08", X"3e", X"78", X"58",
		X"45", X"16", X"93", X"d4", X"df", X"b9", X"1c", X"00", X"06", X"09", X"1b", X"0e", X"2d", X"69", X"89",
		X"70", X"4c", X"28", X"23", X"09", X"07", X"01", X"00", X"07", X"24", X"24", X"06", X"10", X"00", X"00",
		X"48", X"5e", X"07", X"14", X"1e", X"1d", X"3d", X"07", X"00", X"04", X"12", X"61", X"92", X"75", X"88",
		X"30", X"25", X"18", X"00", X"2e", X"72", X"63", X"32", X"2a", X"28", X"79", X"0c", X"61", X"93", X"70",
		X"4d", X"b1", X"b2", X"3c", X"72", X"cd", X"72", X"c6", X"94", X"78", X"5b", X"05", X"be", X"c4", X"67",
		X"9f", X"59", X"a4", X"41", X"00", X"2e", X"6f", X"52", X"19", X"36", X"69", X"0d", X"92", X"52", X"82",
		X"1b", X"00", X"00", X"bd", X"e0", X"bf", X"1b", X"00", X"06", X"4c", X"3a", X"03", X"2b", X"4d", X"96",
		X"9f", X"a1", X"80", X"45", X"01", X"0c", X"00", X"00", X"02", X"16", X"26", X"12", X"08", X"00", X"00",
		X"31", X"09", X"36", X"00", X"0a", X"22", X"25", X"1d", X"00", X"00", X"00", X"7e", X"c6", X"5a", X"57",
		X"00", X"32", X"00", X"0f", X"2d", X"3f", X"3d", X"23", X"4f", X"00", X"00", X"00", X"0b", X"43", X"30",
		X"1e", X"b2", X"b1", X"90", X"92", X"d9", X"ee", X"d0", X"b8", X"9b", X"69", X"46", X"ce", X"eb", X"e3",
		X"e5", X"c0", X"ca", X"a5", X"c0", X"04", X"85", X"62", X"09", X"36", X"01", X"64", X"b7", X"63", X"38",
		X"03", X"44", X"66", X"2b", X"a3", X"e6", X"99", X"47", X"13", X"29", X"3c", X"04", X"24", X"4f", X"76",
		X"8f", X"cc", X"ad", X"5a", X"0c", X"04", X"00", X"00", X"0b", X"1e", X"2a", X"05", X"00", X"00", X"00",
		X"50", X"28", X"00", X"0f", X"00", X"00", X"43", X"12", X"12", X"09", X"00", X"7c", X"2a", X"4d", X"44",
		X"01", X"3a", X"00", X"17", X"14", X"0d", X"52", X"00", X"b4", X"60", X"00", X"08", X"04", X"36", X"1e",
		X"11", X"ff", X"c4", X"76", X"d2", X"dd", X"cc", X"e5", X"99", X"62", X"8f", X"fa", X"be", X"6e", X"f2",
		X"ef", X"d7", X"b8", X"66", X"6b", X"86", X"43", X"3e", X"77", X"00", X"05", X"a4", X"80", X"42", X"17",
		X"00", X"19", X"86", X"7f", X"a0", X"ab", X"9c", X"94", X"5a", X"19", X"34", X"32", X"8c", X"8c", X"a9",
		X"83", X"c2", X"d4", X"b6", X"48", X"07", X"00", X"00", X"00", X"0c", X"0f", X"00", X"00", X"00", X"00",
		X"35", X"50", X"00", X"1d", X"26", X"1e", X"35", X"2c", X"26", X"00", X"06", X"04", X"1d", X"36", X"0b",
		X"50", X"50", X"07", X"17", X"11", X"01", X"21", X"28", X"96", X"a2", X"00", X"04", X"00", X"20", X"54",
		X"54", X"5a", X"92", X"a9", X"a8", X"b1", X"80", X"bd", X"b3", X"68", X"00", X"e1", X"e3", X"ea", X"1d",
		X"00", X"c2", X"ec", X"6f", X"53", X"20", X"9a", X"73", X"c4", X"00", X"3b", X"32", X"0e", X"0a", X"46",
		X"0b", X"31", X"28", X"cf", X"e5", X"9a", X"34", X"33", X"2c", X"00", X"11", X"51", X"44", X"72", X"2f",
		X"27", X"96", X"b4", X"af", X"bb", X"3b", X"00", X"00", X"07", X"17", X"26", X"26", X"52", X"00", X"04",
		X"4f", X"63", X"3c", X"00", X"2c", X"79", X"99", X"34", X"1e", X"1f", X"00", X"00", X"4a", X"5f", X"05",
		X"15", X"76", X"33", X"00", X"0c", X"25", X"37", X"0f", X"0a", X"04", X"1f", X"12", X"33", X"42", X"0b",
		X"77", X"a0", X"cc", X"3a", X"fe", X"d2", X"67", X"00", X"00", X"01", X"53", X"37", X"62", X"3f", X"e4",
		X"a0", X"c3", X"3a", X"7e", X"46", X"d9", X"0f", X"62", X"1a", X"5c", X"3b", X"33", X"19", X"2f", X"1f",
		X"5e", X"5e", X"82", X"94", X"73", X"b5", X"d1", X"55", X"4d", X"44", X"00", X"05", X"2c", X"88", X"98",
		X"cf", X"95", X"a0", X"aa", X"97", X"78", X"00", X"06", X"05", X"06", X"3a", X"4f", X"5f", X"00", X"03",
		X"6f", X"55", X"3e", X"83", X"04", X"2d", X"38", X"47", X"1c", X"85", X"62", X"2a", X"2a", X"28", X"0a",
		X"bb", X"f8", X"8d", X"02", X"05", X"2a", X"21", X"76", X"8b", X"44", X"3f", X"33", X"00", X"3c", X"1b",
		X"4a", X"8b", X"a4", X"4c", X"64", X"f6", X"71", X"00", X"00", X"00", X"33", X"6c", X"44", X"3e", X"d5",
		X"c3", X"24", X"aa", X"f8", X"8a", X"84", X"0d", X"02", X"78", X"65", X"3e", X"67", X"35", X"29", X"22",
		X"4a", X"38", X"00", X"5a", X"6e", X"8e", X"c6", X"5a", X"00", X"15", X"2d", X"14", X"00", X"15", X"00",
		X"14", X"10", X"68", X"9e", X"a0", X"54", X"00", X"00", X"00", X"09", X"30", X"58", X"72", X"45", X"3f",
		X"66", X"5d", X"0c", X"7c", X"82", X"1a", X"13", X"04", X"85", X"86", X"87", X"70", X"32", X"59", X"7c",
		X"81", X"d4", X"42", X"07", X"00", X"34", X"61", X"67", X"d9", X"92", X"17", X"78", X"00", X"02", X"5f",
		X"29", X"56", X"20", X"7a", X"26", X"30", X"76", X"00", X"00", X"20", X"10", X"44", X"56", X"8e", X"ef",
		X"00", X"4b", X"c2", X"a3", X"b5", X"56", X"0c", X"42", X"71", X"3b", X"a5", X"30", X"3a", X"18", X"28",
		X"29", X"17", X"1e", X"97", X"52", X"69", X"c2", X"0e", X"c2", X"71", X"2a", X"1d", X"1f", X"0d", X"08",
		X"37", X"42", X"53", X"82", X"ae", X"6c", X"00", X"00", X"00", X"00", X"18", X"44", X"4b", X"38", X"28",
		X"70", X"05", X"21", X"14", X"89", X"9d", X"30", X"2e", X"a7", X"ca", X"a2", X"cd", X"b9", X"9d", X"87",
		X"68", X"a9", X"2b", X"1d", X"10", X"4e", X"74", X"4d", X"5e", X"41", X"0e", X"1d", X"2b", X"1f", X"8a",
		X"0b", X"27", X"30", X"6f", X"62", X"34", X"05", X"22", X"1b", X"48", X"25", X"2a", X"46", X"0c", X"2e",
		X"ad", X"3b", X"0f", X"0e", X"8a", X"0b", X"38", X"72", X"7d", X"78", X"7e", X"49", X"9f", X"0f", X"0e",
		X"16", X"45", X"48", X"6c", X"10", X"38", X"6f", X"38", X"d2", X"b7", X"6e", X"39", X"27", X"00", X"00",
		X"1d", X"26", X"22", X"4e", X"9c", X"a9", X"3e", X"1a", X"00", X"00", X"05", X"19", X"25", X"28", X"2c",
		X"6a", X"00", X"3f", X"48", X"35", X"9d", X"56", X"35", X"00", X"cd", X"f0", X"d9", X"c7", X"fa", X"89",
		X"88", X"97", X"33", X"1e", X"00", X"18", X"30", X"88", X"2a", X"1a", X"00", X"00", X"00", X"1a", X"17",
		X"43", X"17", X"7f", X"9b", X"73", X"14", X"25", X"6e", X"41", X"95", X"56", X"19", X"23", X"47", X"4b",
		X"4b", X"2c", X"62", X"91", X"11", X"2f", X"40", X"80", X"62", X"54", X"65", X"5b", X"00", X"1c", X"02",
		X"32", X"3b", X"3f", X"3a", X"2c", X"0d", X"1b", X"64", X"7d", X"8c", X"79", X"52", X"16", X"00", X"00",
		X"10", X"17", X"17", X"09", X"3f", X"49", X"18", X"0d", X"18", X"2c", X"00", X"00", X"10", X"21", X"37",
		X"84", X"e1", X"3e", X"00", X"1f", X"0e", X"15", X"29", X"49", X"19", X"c9", X"a8", X"92", X"8a", X"fd",
		X"9d", X"b6", X"62", X"6d", X"7b", X"43", X"00", X"5d", X"30", X"17", X"ac", X"90", X"4b", X"07", X"01",
		X"3c", X"d2", X"8c", X"7c", X"21", X"a8", X"db", X"d1", X"c1", X"47", X"14", X"2e", X"51", X"3c", X"5d",
		X"4f", X"1e", X"2d", X"6b", X"b5", X"22", X"58", X"06", X"00", X"67", X"46", X"53", X"15", X"45", X"2b",
		X"21", X"2e", X"4a", X"36", X"4e", X"77", X"47", X"00", X"34", X"71", X"a7", X"25", X"5e", X"75", X"40",
		X"0f", X"1c", X"40", X"68", X"0c", X"0c", X"00", X"01", X"21", X"25", X"01", X"0a", X"1e", X"00", X"00",
		X"4d", X"72", X"a8", X"00", X"57", X"5d", X"00", X"07", X"8a", X"aa", X"b1", X"be", X"35", X"3b", X"46",
		X"d1", X"a3", X"3d", X"25", X"4d", X"50", X"08", X"2d", X"66", X"00", X"43", X"c6", X"b6", X"87", X"00",
		X"93", X"93", X"a3", X"99", X"0c", X"c5", X"d8", X"c3", X"ba", X"68", X"30", X"2c", X"33", X"40", X"56",
		X"91", X"69", X"39", X"11", X"5d", X"15", X"59", X"00", X"3e", X"44", X"3e", X"44", X"14", X"51", X"2e",
		X"0e", X"31", X"0d", X"2e", X"24", X"1e", X"31", X"42", X"0a", X"4a", X"64", X"94", X"c8", X"87", X"52",
		X"36", X"5a", X"99", X"7d", X"7b", X"32", X"00", X"05", X"20", X"0e", X"00", X"00", X"19", X"00", X"00",
		X"56", X"25", X"6c", X"00", X"a6", X"c0", X"bc", X"9a", X"9b", X"8e", X"a2", X"d8", X"69", X"66", X"a6",
		X"ce", X"e4", X"6f", X"56", X"1c", X"24", X"29", X"1a", X"5c", X"29", X"00", X"76", X"cf", X"af", X"b0",
		X"a2", X"56", X"dc", X"3a", X"2d", X"99", X"85", X"ca", X"d7", X"b5", X"0f", X"33", X"28", X"2c", X"22",
		X"45", X"68", X"40", X"59", X"25", X"15", X"2d", X"00", X"33", X"91", X"c0", X"e4", X"20", X"22", X"12",
		X"00", X"00", X"57", X"59", X"45", X"36", X"18", X"00", X"00", X"38", X"8b", X"ad", X"d4", X"c0", X"79",
		X"38", X"5a", X"3a", X"61", X"58", X"3d", X"00", X"23", X"4d", X"2a", X"03", X"00", X"1e", X"00", X"00",
		X"1b", X"0f", X"00", X"00", X"2b", X"9d", X"c8", X"f7", X"e3", X"83", X"54", X"b4", X"fa", X"ff", X"a6",
		X"ec", X"8b", X"37", X"07", X"18", X"12", X"1d", X"09", X"1f", X"33", X"ae", X"a4", X"a4", X"de", X"b7",
		X"d0", X"f2", X"2d", X"17", X"08", X"1a", X"9a", X"a0", X"8b", X"00", X"44", X"06", X"3d", X"23", X"31",
		X"62", X"0e", X"23", X"1d", X"18", X"4e", X"00", X"00", X"52", X"ff", X"c6", X"65", X"70", X"ba", X"a7",
		X"3a", X"41", X"bf", X"8f", X"4d", X"1a", X"28", X"13", X"1c", X"15", X"48", X"c5", X"a4", X"cc", X"e4",
		X"63", X"4e", X"5a", X"36", X"2b", X"11", X"00", X"05", X"4d", X"23", X"0c", X"00", X"0e", X"00", X"00",
		X"30", X"72", X"0d", X"33", X"00", X"0b", X"84", X"c2", X"f4", X"d3", X"be", X"c5", X"e2", X"cd", X"72",
		X"c7", X"c2", X"21", X"20", X"0c", X"11", X"4a", X"2c", X"24", X"8f", X"a9", X"95", X"9f", X"c4", X"78",
		X"a5", X"e7", X"20", X"21", X"17", X"69", X"65", X"80", X"75", X"00", X"41", X"ac", X"7a", X"4f", X"6e",
		X"00", X"00", X"4c", X"20", X"19", X"3f", X"1f", X"99", X"e3", X"24", X"00", X"09", X"43", X"9a", X"61",
		X"df", X"46", X"c0", X"94", X"59", X"00", X"22", X"50", X"1c", X"37", X"51", X"28", X"c2", X"ba", X"c0",
		X"54", X"5e", X"86", X"97", X"79", X"65", X"40", X"4b", X"1b", X"3c", X"0e", X"3c", X"21", X"14", X"00",
		X"68", X"55", X"46", X"69", X"4f", X"8e", X"58", X"d7", X"c4", X"90", X"be", X"f6", X"d9", X"6d", X"7d",
		X"7c", X"f3", X"00", X"25", X"00", X"08", X"2f", X"36", X"37", X"3a", X"40", X"75", X"a5", X"c8", X"cb",
		X"a2", X"fa", X"d4", X"33", X"1b", X"89", X"51", X"47", X"7b", X"26", X"9d", X"73", X"83", X"a3", X"85",
		X"00", X"60", X"84", X"6c", X"24", X"a4", X"ba", X"76", X"12", X"06", X"81", X"b2", X"00", X"c2", X"a0",
		X"97", X"d8", X"94", X"ff", X"a5", X"00", X"1a", X"43", X"66", X"ae", X"ad", X"b4", X"b9", X"cc", X"58",
		X"59", X"db", X"db", X"b0", X"4f", X"24", X"0e", X"10", X"0c", X"25", X"02", X"36", X"35", X"00", X"00",
		X"38", X"14", X"53", X"9b", X"df", X"e1", X"cd", X"9f", X"e7", X"4e", X"99", X"a1", X"dd", X"d7", X"7a",
		X"70", X"9b", X"00", X"33", X"15", X"1f", X"3f", X"14", X"31", X"28", X"04", X"25", X"53", X"86", X"c8",
		X"de", X"d0", X"ee", X"ce", X"0c", X"36", X"cf", X"c1", X"b4", X"ee", X"66", X"54", X"93", X"3d", X"b2",
		X"ca", X"95", X"b8", X"3d", X"21", X"4d", X"23", X"23", X"51", X"73", X"ff", X"55", X"9a", X"b3", X"dc",
		X"e3", X"f9", X"dd", X"ff", X"5e", X"00", X"0d", X"42", X"91", X"c1", X"c1", X"d6", X"ef", X"ce", X"44",
		X"0b", X"be", X"cc", X"c4", X"c4", X"98", X"2f", X"00", X"26", X"1f", X"00", X"00", X"1e", X"00", X"00",
		X"38", X"00", X"af", X"7b", X"ca", X"d9", X"e9", X"d5", X"ce", X"00", X"81", X"fc", X"bc", X"df", X"de",
		X"31", X"16", X"00", X"00", X"05", X"00", X"29", X"65", X"2f", X"33", X"00", X"60", X"3f", X"7b", X"88",
		X"ef", X"d6", X"b8", X"b8", X"52", X"14", X"ff", X"df", X"ed", X"ff", X"be", X"9a", X"9c", X"61", X"35",
		X"f1", X"e7", X"ec", X"0e", X"3e", X"23", X"53", X"80", X"5b", X"51", X"ee", X"7e", X"2f", X"76", X"66",
		X"ca", X"f6", X"15", X"7f", X"6c", X"00", X"63", X"96", X"5c", X"5d", X"76", X"9b", X"53", X"43", X"f1",
		X"90", X"d4", X"d6", X"a2", X"19", X"10", X"00", X"00", X"16", X"1e", X"00", X"00", X"08", X"00", X"00",
		X"32", X"24", X"76", X"6f", X"64", X"ef", X"ff", X"a3", X"91", X"af", X"dd", X"c1", X"fb", X"d2", X"b0",
		X"00", X"00", X"04", X"05", X"00", X"0e", X"38", X"56", X"2e", X"16", X"26", X"a5", X"47", X"9c", X"75",
		X"a7", X"b7", X"a2", X"07", X"97", X"8d", X"c9", X"e9", X"58", X"a6", X"ff", X"ca", X"96", X"96", X"f9",
		X"be", X"e9", X"e7", X"00", X"4c", X"75", X"6a", X"37", X"9b", X"f1", X"be", X"94", X"58", X"55", X"d2",
		X"47", X"c4", X"14", X"e7", X"e1", X"3d", X"2a", X"5d", X"4a", X"65", X"57", X"7f", X"27", X"00", X"b5",
		X"8d", X"c7", X"c2", X"ff", X"3b", X"00", X"00", X"00", X"36", X"1f", X"00", X"00", X"00", X"30", X"5f",
		X"1c", X"61", X"5c", X"72", X"82", X"bc", X"29", X"ad", X"b6", X"9d", X"95", X"cb", X"cb", X"d4", X"14",
		X"29", X"05", X"02", X"17", X"16", X"0d", X"28", X"00", X"2d", X"07", X"88", X"a7", X"b8", X"5f", X"40",
		X"79", X"88", X"a4", X"c9", X"cd", X"b2", X"ed", X"b1", X"54", X"1b", X"b9", X"d6", X"84", X"6d", X"93",
		X"bc", X"b8", X"f6", X"8b", X"25", X"35", X"0a", X"b1", X"7b", X"c7", X"e1", X"77", X"ab", X"53", X"45",
		X"49", X"be", X"f4", X"c0", X"c4", X"5a", X"19", X"0f", X"3a", X"6c", X"7f", X"2c", X"37", X"50", X"b5",
		X"a4", X"98", X"60", X"a0", X"e9", X"24", X"00", X"00", X"20", X"00", X"00", X"00", X"00", X"56", X"53",
		X"6c", X"66", X"41", X"4a", X"20", X"2e", X"39", X"b8", X"c2", X"d9", X"a8", X"c9", X"91", X"b0", X"2c",
		X"1e", X"06", X"1a", X"28", X"25", X"18", X"13", X"1d", X"11", X"11", X"20", X"3e", X"00", X"25", X"48",
		X"53", X"7b", X"2d", X"9d", X"b6", X"bb", X"b3", X"ce", X"6f", X"e6", X"c2", X"da", X"99", X"7d", X"a4",
		X"66", X"3a", X"e4", X"f2", X"35", X"00", X"24", X"53", X"6f", X"ff", X"d0", X"3d", X"00", X"07", X"00",
		X"4a", X"a0", X"b7", X"e7", X"a3", X"4f", X"4d", X"50", X"50", X"70", X"41", X"00", X"66", X"00", X"69",
		X"d0", X"22", X"06", X"35", X"b3", X"5e", X"48", X"2b", X"16", X"03", X"0c", X"1b", X"09", X"42", X"3b",
		X"1b", X"22", X"25", X"5d", X"60", X"32", X"17", X"28", X"ba", X"c2", X"43", X"56", X"e2", X"9d", X"74",
		X"2c", X"21", X"0d", X"00", X"12", X"00", X"06", X"0b", X"00", X"1b", X"03", X"00", X"20", X"29", X"0e",
		X"04", X"00", X"4b", X"65", X"b9", X"a2", X"a6", X"a1", X"ff", X"d7", X"8a", X"86", X"76", X"63", X"22",
		X"36", X"3a", X"50", X"ff", X"96", X"0a", X"3e", X"44", X"00", X"e4", X"00", X"39", X"2f", X"0d", X"20",
		X"27", X"6f", X"85", X"ce", X"26", X"40", X"45", X"6c", X"89", X"2f", X"00", X"2b", X"00", X"0e", X"1e",
		X"53", X"05", X"02", X"16", X"5d", X"be", X"0f", X"12", X"09", X"0f", X"00", X"00", X"00", X"3b", X"37",
		X"30", X"1b", X"0c", X"54", X"73", X"12", X"0f", X"00", X"0f", X"a6", X"29", X"56", X"36", X"d1", X"6e",
		X"30", X"00", X"03", X"09", X"11", X"00", X"00", X"14", X"00", X"1f", X"09", X"0f", X"29", X"19", X"08",
		X"19", X"30", X"00", X"00", X"fa", X"e3", X"c3", X"ec", X"a0", X"ff", X"98", X"7d", X"4f", X"02", X"0f",
		X"ff", X"d6", X"29", X"e6", X"1e", X"33", X"58", X"45", X"03", X"00", X"0f", X"5b", X"25", X"1c", X"54",
		X"2d", X"5c", X"68", X"ac", X"00", X"38", X"49", X"95", X"75", X"00", X"67", X"27", X"00", X"1d", X"2a",
		X"0c", X"05", X"10", X"1d", X"00", X"4d", X"00", X"16", X"20", X"10", X"00", X"04", X"05", X"52", X"69",
		X"4f", X"00", X"00", X"00", X"5a", X"63", X"1c", X"0d", X"56", X"6d", X"43", X"15", X"c6", X"b1", X"a2",
		X"66", X"00", X"02", X"17", X"05", X"04", X"03", X"0f", X"12", X"1e", X"02", X"00", X"35", X"47", X"00",
		X"14", X"46", X"14", X"29", X"e5", X"d5", X"ff", X"df", X"63", X"ff", X"d5", X"b2", X"74", X"05", X"ab",
		X"c2", X"aa", X"28", X"70", X"44", X"31", X"7a", X"36", X"2f", X"00", X"1b", X"31", X"2e", X"23", X"32",
		X"37", X"3b", X"38", X"42", X"00", X"2b", X"77", X"74", X"00", X"42", X"52", X"00", X"05", X"18", X"12",
		X"18", X"00", X"00", X"00", X"52", X"00", X"57", X"03", X"08", X"00", X"00", X"00", X"0b", X"60", X"67",
		X"17", X"0e", X"05", X"06", X"01", X"48", X"03", X"0a", X"49", X"4e", X"61", X"8c", X"da", X"e0", X"60",
		X"6b", X"53", X"00", X"00", X"04", X"00", X"13", X"13", X"0e", X"0e", X"05", X"00", X"35", X"00", X"0b",
		X"27", X"0b", X"20", X"0b", X"40", X"ac", X"5d", X"2c", X"10", X"73", X"cb", X"b3", X"3e", X"13", X"b9",
		X"a2", X"d1", X"ff", X"7e", X"da", X"8f", X"86", X"8c", X"e0", X"4e", X"00", X"33", X"2e", X"1a", X"6a",
		X"76", X"1a", X"27", X"80", X"00", X"45", X"46", X"00", X"54", X"28", X"09", X"20", X"00", X"00", X"00",
		X"1f", X"c4", X"89", X"91", X"11", X"3b", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5a", X"52",
		X"15", X"0a", X"13", X"0e", X"08", X"2a", X"14", X"27", X"4b", X"4f", X"51", X"1f", X"5b", X"bf", X"7d",
		X"76", X"10", X"0e", X"00", X"04", X"18", X"0c", X"00", X"19", X"00", X"70", X"b1", X"62", X"b0", X"1f",
		X"0b", X"43", X"2c", X"18", X"00", X"55", X"29", X"ef", X"42", X"22", X"04", X"8c", X"93", X"a6", X"b5",
		X"c3", X"b7", X"6f", X"78", X"60", X"dc", X"a8", X"55", X"92", X"c5", X"00", X"31", X"1f", X"5c", X"a8",
		X"40", X"30", X"3f", X"21", X"05", X"23", X"04", X"1d", X"55", X"31", X"00", X"00", X"00", X"05", X"0c",
		X"5d", X"39", X"0a", X"00", X"0f", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"50", X"55",
		X"00", X"00", X"00", X"13", X"28", X"1d", X"2c", X"16", X"19", X"11", X"5b", X"4e", X"63", X"17", X"4f",
		X"6c", X"62", X"00", X"06", X"00", X"00", X"40", X"11", X"13", X"14", X"b5", X"1e", X"c6", X"f4", X"ff",
		X"00", X"1b", X"2b", X"1b", X"6a", X"10", X"21", X"d4", X"ff", X"3f", X"23", X"5d", X"e6", X"77", X"bc",
		X"f0", X"b4", X"b6", X"85", X"c3", X"d6", X"5b", X"48", X"c1", X"b7", X"d4", X"ce", X"a5", X"0b", X"45",
		X"44", X"1d", X"49", X"34", X"42", X"00", X"16", X"1b", X"28", X"61", X"6f", X"68", X"69", X"0f", X"15",
		X"00", X"11", X"48", X"3b", X"35", X"16", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"33", X"27",
		X"00", X"00", X"00", X"15", X"2e", X"0b", X"19", X"1f", X"12", X"08", X"9f", X"45", X"6f", X"3d", X"a4",
		X"6c", X"00", X"00", X"02", X"0c", X"13", X"4f", X"00", X"09", X"2b", X"a9", X"c7", X"65", X"d4", X"ff",
		X"ed", X"09", X"0f", X"67", X"54", X"0c", X"16", X"3a", X"b4", X"13", X"13", X"98", X"84", X"62", X"4e",
		X"e4", X"cf", X"e0", X"bb", X"c8", X"d1", X"93", X"10", X"c2", X"bb", X"ff", X"df", X"f1", X"3b", X"2d",
		X"2b", X"15", X"25", X"2a", X"38", X"30", X"2b", X"00", X"01", X"20", X"15", X"21", X"6e", X"56", X"3e",
		X"39", X"09", X"1a", X"0d", X"10", X"00", X"26", X"25", X"10", X"00", X"00", X"00", X"00", X"22", X"23",
		X"5a", X"00", X"00", X"00", X"1c", X"00", X"00", X"28", X"00", X"00", X"6d", X"59", X"24", X"00", X"00",
		X"1f", X"00", X"00", X"00", X"12", X"4c", X"38", X"00", X"0a", X"17", X"17", X"f3", X"ef", X"bd", X"9e",
		X"e6", X"e3", X"a5", X"e0", X"bf", X"04", X"4b", X"ac", X"10", X"26", X"8d", X"12", X"d2", X"ec", X"3b",
		X"de", X"cf", X"b6", X"d7", X"d3", X"a1", X"bc", X"56", X"d9", X"e8", X"d7", X"e8", X"c8", X"74", X"00",
		X"32", X"11", X"20", X"59", X"40", X"2a", X"17", X"00", X"00", X"00", X"01", X"01", X"36", X"00", X"0c",
		X"0a", X"28", X"39", X"10", X"00", X"37", X"35", X"3d", X"36", X"38", X"12", X"0e", X"10", X"12", X"09",
		X"5a", X"3b"
	);

	signal clock_counter      : natural := 0;
	signal clock_counter_stop : natural := 0;

	signal errors_nb : natural := 0;

	-- Defined in VHDL 2008, not handled by GHDL
	function to_string(sv: std_logic_vector) return string is
		variable bv: bit_vector(sv'range) := to_bitvector(sv);
		variable lp: line;
	begin
		write(lp, bv);
		return lp.all;
	end;

begin

	-- Instantiation of the main component
	top_i : top port map (
		-- Access 'clock' model 'clock'
		clock => clock,
		-- Access 'reset' model 'reset'
		reset => reset,
		-- Access 'start' model 'start'
		start => start,
		-- Access 'stdin' model 'fifo_in'
		stdin_data => stdin_data,
		stdin_rdy => stdin_rdy,
		stdin_ack => stdin_ack,
		-- Access 'stdout' model 'fifo_out'
		stdout_data => stdout_data,
		stdout_rdy => stdout_rdy,
		stdout_ack => stdout_ack
	);

	-- Functionality for top-level access 'clock' model 'clock'
	-- Generation of clock: 100MHz (note: arbitrary value)
	clock <= clock_next after 5 ns;
	clock_next <= not clock when clock_counter_stop = 0 or clock_counter <= clock_counter_stop else '0';

	-- Clock counter and global messages
	process (clock)
		-- To print simulation messages
		variable l : line;
	begin

		-- Increment clock counter
		if rising_edge(clock) then

			clock_counter <= clock_counter + 1;

			if simu_disp_cycles = '1' then
				-- Write simulation message
				write(l, string'("INFO clock cycle "));
				write(l, clock_counter);
				writeline(output, l);
			end if;

		end if;

		-- Messages
		if falling_edge(clock) then

			if clock_counter > simu_max_cycles then
				report "ERROR Too many cycles simulated. Stopping simulation." severity failure;
			end if;

			if clock_counter < reset_cycles then
				report "INFO Reset" severity note;
			end if;

			if clock_counter = reset_cycles then
				report "INFO Start" severity note;
			end if;

		end if;

	end process;

	-- Functionality for top-level access 'reset' model 'reset'
	-- Generation of reset
	reset <= '1' when clock_counter < reset_cycles else '0';

	-- Functionality for top-level access 'start' model 'start'
	-- Generation of start
	start <= '1';

	-- Functionality for top-level access 'stdin' model 'fifo_in'
	-- FIFO stdin
	-- Sending inputs

	stdin_vector <= stdin_vectors(stdin_vector_idx) when stdin_vector_idx < stdin_vectors_nb else (others => '0');
	stdin_data <= stdin_vector(7 downto 0);

	stdin_ack <= '1' when reset = '0' and stdin_vector_idx < stdin_vectors_nb else '0';

	process (clock)
		-- To print simulation messages
		variable l : line;
	begin

		if rising_edge(clock) then

			if stdin_vector_idx < stdin_vectors_nb then

				if stdin_rdy = '1' and stdin_ack = '1' and reset = '0' then

					-- Write simulation message
					write(l, string'("INFO Input vector "));
					write(l, stdin_vector_idx);
					write(l, string'(" at cycle "));
					write(l, clock_counter);
					writeline(output, l);

					if stdin_vector_idx = 0 then
						write(l, string'("INFO First input vector sent at clock cycle "));
						write(l, clock_counter);
						writeline(output, l);
					end if;

					if stdin_vector_idx = stdin_vectors_nb - 1 then
						write(l, string'("INFO Last input vector sent at clock cycle "));
						write(l, clock_counter);
						writeline(output, l);
					end if;

					-- Increase vector index
					stdin_vector_idx <= stdin_vector_idx + 1;

				end if;  -- Handshake

			else

				if stdin_rdy = '1' and reset = '0' then
					if simu_err_end_in = '1' then
						report "ERROR Out of input vectors. Stopping simulation." severity failure;
					end if;
				end if;  -- Handshake

			end if;

		end if;

	end process;

	-- Functionality for top-level access 'stdout' model 'fifo_out'
	-- FIFO stdout
	-- Checking outputs

	-- Always enable output FIFO
	stdout_ack <= '1' when stdout_vector_idx < stdout_vectors_nb and reset = '0' else '0';

	stdout_vector <= stdout_vectors(stdout_vector_idx) when stdout_vector_idx < stdout_vectors_nb else (others => '0');

	-- Check outputs
	process (clock)
		variable l : line;
	begin

		if rising_edge(clock) then

			if stdout_vector_idx < stdout_vectors_nb then

				if stdout_rdy = '1' and stdout_ack = '1' and reset = '0' then

					if stdout_data = stdout_vector(7 downto 0) then
						-- The vector is verified

						write(l, string'("INFO Output nb "));
						write(l, stdout_vector_idx);
						write(l, string'(" at cycle "));
						write(l, clock_counter);
						write(l, string'(" (check OK)"));
						write(l, string'(" Obtained "));
						write(l, to_string(stdout_data));
						writeline(output, l);

					else
						-- An error is detected

						write(l, string'("ERROR Output nb "));
						write(l, stdout_vector_idx);
						write(l, string'(" at cycle "));
						write(l, clock_counter);
						writeline(output, l);

						write(l, string'("  Obtained "));
						write(l, to_string(stdout_data));
						writeline(output, l);
						write(l, string'("  Expected "));
						write(l, to_string(stdout_vector(7 downto 0)));
						writeline(output, l);

						errors_nb <= errors_nb + 1;

						--report "ERROR A simulation error was found." severity failure;

					end if;

					if stdout_vector_idx = stdout_vectors_nb - 1 then

						write(l, string'("INFO Last output vector read at cycle "));
						write(l, clock_counter);
						writeline(output, l);

						report "INFO Stopping simulation." severity note;

						clock_counter_stop <= clock_counter + 3;

					end if;

					-- Increase vector index
					stdout_vector_idx <= stdout_vector_idx + 1;

				end if;  -- FIFO handshake

			else
				-- All vectors have been read

				if errors_nb > 0 then
					write(l, string'("ERROR Number of errors found : "));
					write(l, errors_nb);
					writeline(output, l);
					report "ERROR Simulation errors were found." severity failure;
				end if;

			end if;  -- Check all vectors read

		end if;  -- Clock

	end process;

end augh;

