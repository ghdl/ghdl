﻿-- This is utf-8 encoding, with a BOM.

package p1 is
end p1;

