architecture;s';