package p is
  function B return p'xx;
end;

