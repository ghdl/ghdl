
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc43.vhd,v 1.2 2001-10-26 16:29:54 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c04s03b01x01p02n01i00043ent IS
END c04s03b01x01p02n01i00043ent;

ARCHITECTURE c04s03b01x01p02n01i00043arch OF c04s03b01x01p02n01i00043ent IS
  -- constant integer:integer := 1;  -- No_failure_here
  -- According to scopes and visibility rules, this test is not correct.
  constant integer:natural := 1;
BEGIN
  TESTING: PROCESS
  BEGIN
    assert NOT(integer = 1)
      report "***PASSED TEST: c04s03b01x01p02n01i00043" 
      severity NOTE;
    assert (integer = 1)
      report "***FAILED TEST:c04s03b01x01p02n01i00043 - Constant declaration test failed."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c04s03b01x01p02n01i00043arch;
