package Util is
  type integer_list_t is array (natural range <>) of integer;
end package;
