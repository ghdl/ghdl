entity test_val is end test_val; 
architecture test of test_val is 
signal t : time := time'value("123 fs"); 
begin 
end test; 
