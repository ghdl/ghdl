--library osvvm;
use work.ResolutionPkg.all;

entity Resolution_TB is
end Resolution_TB;

architecture none of Resolution_TB is
begin
end none;
