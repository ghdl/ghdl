entity e is end;

architecture a of e is
begin
end;

