architecture arch of ent is
  signal s1 : bit;  --  comment for :s1:
  --  Also for :s1:
  signal s2: natural;
begin
end arch;
