
-- Copyright (C) 2002 Morgan Kaufmann Publishers, Inc

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

entity tb_full_adder is
end entity tb_full_adder;


library util;  use util.stimulus_generators.all;

architecture test of tb_full_adder is

  signal a, b, c_in, s, c_out : bit;
  signal test_vector : bit_vector(1 to 3);

begin

  dut : entity work.full_adder
    port map ( a => a, b => b, c_in => c_in, s => s, c_out => c_out );

  all_possible_values ( test_vector, 10 ns );

  (a, b, c_in) <= test_vector;

end architecture test;
