-- Author:  Patrick Lehmann
-- License: MIT
--
-- undocumented
--
context StopWatch_ctx is
	library lib_Utilities;
	context lib_Utilities.Utilities_ctx;

	use work.StopWatch_pkg.all;
end context;
