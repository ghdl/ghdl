use work.MemorySupportPkg.all;

entity ent is
end;

architecture behav of ent is
  constant c : MemBlockType := InitMemoryBaseType_X (3, 2);
begin
end;
