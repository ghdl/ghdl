
-- Copyright (C) 1996 Morgan Kaufmann Publishers, Inc

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: ch_04_ch_04_04.vhd,v 1.2 2001-10-26 16:29:33 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

entity ch_04_04 is

end entity ch_04_04;


----------------------------------------------------------------


architecture test of ch_04_04 is
begin


  process_04_1_i : process is

                             -- code from book:

                             type A is array (1 to 4, 31 downto 0) of boolean;

                           -- end of code from book

                           variable free_map : bit_vector(1 to 10) := "0011010110";
                           variable count : natural;

  begin

    -- code from book (just the conditions):

    assert A'left(1) = 1;      assert A'low(1) = 1;
    assert A'right(2) = 0 ;    assert A'high(2) = 31;

    assert A'length(1) = 4;    assert A'length(2) = 32;

    assert A'ascending(1) = true;    assert A'ascending(2) = false;

    assert A'low = 1;    assert A'length = 4;

    --

    count := 0;
    for index in free_map'range loop
      if free_map(index) = '1' then
        count := count + 1;
      end if;
    end loop;

    -- end of code from book

    wait;
  end process process_04_1_i;


end architecture test;
