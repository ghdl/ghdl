
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1442.vhd,v 1.2 2001-10-26 16:29:41 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c08s07b00x00p02n01i01442ent IS
END c08s07b00x00p02n01i01442ent;

ARCHITECTURE c08s07b00x00p02n01i01442arch OF c08s07b00x00p02n01i01442ent IS

begin
  TESTING: process
    variable k : integer := 0;
    variable m : integer := 6;
    variable j : boolean := TRUE;
  begin
    if m > 5 then
      case j is
        when TRUE   => k := 1;
        when FALSE   => NULL;
      end case;
    end if;
    assert NOT(k = 1)
      report "***PASSED TEST: c08s07b00x00p02n01i01442"
      severity NOTE;
    assert (k = 1)
      report "***FAILED TEST: c08s07b00x00p02n01i01442 - CASE statement to be sequence statements of IF statement" 
      severity ERROR;
    wait;
  end process TESTING;

END c08s07b00x00p02n01i01442arch;
