package p is
  function log2(
    -- :param1: we also want to document parameters too
    param1 : integer;
    param2 : boolean
    ) return natural;
end p;


