
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc344.vhd,v 1.2 2001-10-26 16:29:53 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s02b01x00p09n01i00344ent IS
END c03s02b01x00p09n01i00344ent;

ARCHITECTURE c03s02b01x00p09n01i00344arch OF c03s02b01x00p09n01i00344ent IS

BEGIN
  TESTING: PROCESS
    type       T_A1_S       is ARRAY(INTEGER range <>) of INTEGER;
    subtype    ST_A1_S    is T_A1_S(INTEGER range 1 to 3);

    variable    V_A1_S       : ST_A1_S;
  BEGIN
    V_A1_S(1) := 11;
    V_A1_S(2) := 22;
    V_A1_S(3) := 33;
    wait for 5 ns;
    assert NOT(   V_A1_S(1) = 11   and
                  V_A1_S(2) = 22   and
                  V_A1_S(3) = 33   )
      report "***PASSED TEST: c03s02b01x00p09n01i00344"
      severity NOTE;
    assert (   V_A1_S(1) = 11   and
               V_A1_S(2) = 22   and
               V_A1_S(3) = 33   )
      report "***FAILED TEST: c03s02b01x00p09n01i00344 - For each possible index value there should be a distinct element."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s02b01x00p09n01i00344arch;
