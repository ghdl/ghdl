entity g is
  generic(type stream0t);
  port(t:t stream0t);
end;

architecture t of g is
  type e is array(0)of m;
  signal w:r range 0 to 0;
  signal r:r range 0 to 0;
  signal m:n;
begin
  y(0);
  process(a)
  begin
    if(0)then
      if 0 then(0)<=0;
      end if;
    end if;
  end process;
end;
