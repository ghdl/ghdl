package aa2 is
constant a : bit_vector(0 to 1) := ('0', '1');
constant b : bit_vector(0 to 0) := a(integer range 0 to 0);
end package aa2;
