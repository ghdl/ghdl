package p is
  --  Comment for the decl.
  constant c1 : natural := 3;
end p;
