entity hello is
  error;
end hello;
