library ieee;
use ieee.std_logic_unsigned;

entity tb is
end tb;
