package function begin c';