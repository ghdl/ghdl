library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ent is
    port (
    aaa : in std_logic);
end ent;

architecture structure of ent is
begin
end structure;
