
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2642.vhd,v 1.2 2001-10-26 16:29:49 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

entity THIS_IS_A_PRETTY_LONG_NAME_FOR_AN_ENTI is
end;

entity THIS_IS_A_PRETTY_LONG_NAME_FOR_AN_ENTIT is
end;

entity THIS_IS_A_PRETTY_LONG_NAME_FOR_AN_ENTITY is
end;

entity This_Entity_Name_Is_Not_Long is
end;

architecture This_Arch_Name_Is_Not_Long of This_Entity_Name_Is_Not_Long is
begin
end;

ENTITY c13s03b01x00p02n01i02642ent IS
END c13s03b01x00p02n01i02642ent;

ARCHITECTURE c13s03b01x00p02n01i02642arch OF c13s03b01x00p02n01i02642ent IS

BEGIN
  TESTING: PROCESS
  BEGIN
    assert FALSE 
      report "***PASSED TEST: c13s03b01x00p02n01i02642" 
      severity NOTE;
    wait;
  END PROCESS TESTING;

END c13s03b01x00p02n01i02642arch;
