entity e is
end entity;

architecture a of e is
begin
  end: std.env.stop;
end architecture;

package p is
end package;
