
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1074.vhd,v 1.2 2001-10-26 16:30:29 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c06s04b00x00p03n04i01074ent IS
END c06s04b00x00p03n04i01074ent;

ARCHITECTURE c06s04b00x00p03n04i01074arch OF c06s04b00x00p03n04i01074ent IS
BEGIN
  TESTING: PROCESS
    constant C1 : STRING    := "ABCDEFGH";
    variable V1 : CHARACTER;
    variable q  : integer    := 9;
  BEGIN
    V1 := C1(1);
    assert V1 = 'A' 
      report "FAIL: first index";
    V1 := C1(q);                    -- should result in index error
    assert FALSE 
      report "***FAILED TEST: c06s04b00x00p03n04i01074- Index value should belong to the range of the corresponding index range of the array." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c06s04b00x00p03n04i01074arch;
