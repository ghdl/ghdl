
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc503.vhd,v 1.2 2001-10-26 16:29:55 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s02b02x00p03n01i00503ent IS
END c03s02b02x00p03n01i00503ent;

ARCHITECTURE c03s02b02x00p03n01i00503arch OF c03s02b02x00p03n01i00503ent IS
  type R2 is record
               R11,R12 : INTEGER;
               R21,R22,R23 : BOOLEAN;
             end record;
BEGIN
  TESTING: PROCESS
    variable k : R2;
  BEGIN
    k.R11   := 1;
    k.R12   := 2;
    k.R21   := true;
    k.R22   := false;
    k.R23   := true;
    wait for 2 ns;
    assert NOT(k.R11=1 and k.R12=2 and k.R21=true and k.R22=false and k.R23=true)
      report "***PASSED TEST: c03s02b02x00p03n01i00503"
      severity NOTE;
    assert (k.R11=1 and k.R12=2 and k.R21=true and k.R22=false and k.R23=true)
      report "***FAILED TEST: c03s02b02x00p03n01i00503 - A multiple object declaration is equivalent to a sequence of the corresponding number of single object declarations."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s02b02x00p03n01i00503arch;
