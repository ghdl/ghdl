architecture function(0is;0package