
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc1732.vhd,v 1.2 2001-10-26 16:29:43 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c09s03b00x00p14n01i01732ent IS
END c09s03b00x00p14n01i01732ent;

ARCHITECTURE c09s03b00x00p14n01i01732arch OF c09s03b00x00p14n01i01732ent IS
  signal    s1 : bit;
  signal    s2 : integer;
  signal    s3 : integer;

  procedure unguarded_proc (where : in integer; signal here : out integer) is
  begin
    if where = 1 then
      here <= 5;
    else
      here <= 6;
    end if;
  end;

BEGIN
  s3   <= 1 after 20 ns;

  block_label1 : BLOCK ( s1 = '1' )
  begin
    unguarded_proc (s3,s2);
  end block block_label1;

  TESTING: PROCESS(s2)
  BEGIN
    if (now > 1 ns) then
      assert NOT( s2=5 )
        report "***PASSED TEST: c09s03b00x00p14n01i01732"
        severity NOTE;
      assert ( s2=5 )
        report "***FAILED TEST: c09s03b00x00p14n01i01732 - The value of an implicitly declared signal GUARD has no effect on evaluation of a concurrent procedure call."
        severity ERROR;
    end if;
  END PROCESS TESTING;

END c09s03b00x00p14n01i01732arch;
