library ieee;use ieee.std_logic_1164;entity d is
port(s:std'r);end entity;architecture c of t is
begin
t;end architecture;