package std_logic_textio is
  -- empty.
end std_logic_textio;
