entity e is
end;

architecture behav of e is
begin
  assert g[](0);
end;
