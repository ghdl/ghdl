context work.prj;

entity ent1 is
end ent1;

architecture behav of ent1 is
  signal s : std_ulogic;
begin
end behav;
