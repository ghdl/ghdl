library ieee;
use ieee.all.common.workall;
entity icache is end;
