package n is
  generic(package g is new n generic map(<>));
  function t return l;
end;
