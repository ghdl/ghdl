entity tb is
end tb;

architecture behavioral of tb is
   subtype int30 is integer range -1 to 0**0;
begin
 end behavioral;

