
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc3162.vhd,v 1.2 2001-10-26 16:29:52 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c14s01b00x00p07n01i03162ent IS
END c14s01b00x00p07n01i03162ent;

ARCHITECTURE c14s01b00x00p07n01i03162arch OF c14s01b00x00p07n01i03162ent IS

BEGIN
  TESTING: PROCESS

    subtype BTRUE    is BOOLEAN range TRUE to TRUE;
    subtype ST    is INTEGER range -5 to 20;

    type E is (A,B,C,D);
    type P is range 1 to 24
      units
        U;
        X=3 U;
        Y=2 X;
      end units;

  BEGIN
    wait for 5 ns;
    assert NOT(       (E'BASE'LEFT   =E'LEFT)
                      and    (REAL'BASE'HIGH   =REAL'HIGH)
                      and    (E'BASE'POS(C)   =E'POS(C))
                      and    (ST'BASE'VAL(1)   =INTEGER'VAL(1))
                      and    (INTEGER'BASE'PRED(1)   =INTEGER'PRED(1))
                      and    (P'BASE'SUCC(2 Y)   =P'SUCC(2 Y)))
      report "***PASSED TEST: /src/ch14/sc01/p007/s010101.vhd"
      severity NOTE;
    assert (       (E'BASE'LEFT   =E'LEFT)
                   and    (REAL'BASE'HIGH   =REAL'HIGH)
                   and    (E'BASE'POS(C)   =E'POS(C))
                   and    (ST'BASE'VAL(1)   =INTEGER'VAL(1))
                   and    (INTEGER'BASE'PRED(1)   =INTEGER'PRED(1))
                   and    (P'BASE'SUCC(2 Y)   =P'SUCC(2 Y)))
      report "***FAILED TEST: c14s01b00x00p07n01i03162 - Result of T'BASE must be same as the base type of T."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c14s01b00x00p07n01i03162arch;
