architecture	if''h';