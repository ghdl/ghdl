library ieee;use ieee.std_logic_1164.all;entity dut is
port(sig_i:std_logic_vector;sig_o:out std_logic_vector);end entity;architecture a of dut is
begin	sig_o<=sig_i;end architecture;library ieee;use ieee.std_logic_1164;entity tb is
end entity;architecture h of tb is
signal n:std'r(0);signal s:s(0);begin process	begin
end process;t(0);end architecture;