-- This is standard 7bit ascii encoding

package p1 is
end p1;
