package p is

  constant c : natural := 1;

  --  Comment
  type vec is array(natural range <>) of bit_vector(0 to 1);
end p;
