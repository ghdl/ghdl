entity reserved3 is
end;

architecture behav of reserved3 is
  signal protected : bit;
begin
  process
  begin
    wait;
  end process;
end behav;
