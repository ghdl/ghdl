
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2399.vhd,v 1.2 2001-10-26 16:29:47 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c07s03b02x00p08n01i02399ent IS
END c07s03b02x00p08n01i02399ent;

ARCHITECTURE c07s03b02x00p08n01i02399arch OF c07s03b02x00p08n01i02399ent IS

BEGIN
  TESTING: PROCESS
    type rec is record
                  ele_2 : real;
                  ele_3 : boolean;
                end record;
    variable v23 : rec;
  BEGIN
    v23 := (ele_2 => 2.3, ele_3 => True); -- No_failure_here
    assert NOT((v23.ele_2=2.3) and (v23.ele_3=TRUE)) 
      report "***PASSED TEST: c07s03b02x00p08n01i02399" 
      severity NOTE;
    assert ((v23.ele_2=2.3) and (v23.ele_3=TRUE)) 
      report "***FAILED TEST: c07s03b02x00p08n01i02399 - Element associations by an element simple name is allowed only in record aggregates."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c07s03b02x00p08n01i02399arch;
