package mypkg is
	type foo;
	type foo_acc is access foo;

	type foo is protected
	end protected;
end package mypkg;
