package p is
  type state_t is
    (
      --  Comment for :s1:
      s1,
      s2,
      s3);
end p;
