architecture�0for(4000000000x"