entity repro3 is
end;

architecture behav of repro3 is
begin
   process
   begin
    "and" (true, false);
   end process;
end;
