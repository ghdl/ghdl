
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2891.vhd,v 1.2 2001-10-26 16:30:23 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c02s01b01x00p05n01i02891ent IS
  PORT ( d  : IN  bit;
         q  : OUT bit);
END c02s01b01x00p05n01i02891ent;

ARCHITECTURE c02s01b01x00p05n01i02891arch OF c02s01b01x00p05n01i02891ent IS
  function func1 (signal p1 : in bit) return bit;
  function func2 (signal p1 : buffer bit) return bit;

  function func1 (signal p1 : in bit) return bit is
    variable v1 : bit;
  begin
    v1 := p1;
    return (v1);
  end;

  function func2 (signal p1 : buffer bit) return bit is
    variable v1 : bit;
  begin
    v1 := p1;
    return (v1);
  end;
BEGIN
  func1 (d);
  func2 (d);
  q <= d;

  TESTING: PROCESS
  BEGIN
    assert FALSE
      report "***FAILED TEST: c02s01b01x00p05n01i02891 - Buffer is not an allowed mode for formal parameters of a function."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c02s01b01x00p05n01i02891arch;
