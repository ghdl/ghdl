library ieee;
use ieee.std_logic_1164.all;

package apkg is

    component acomp is
        port (x: in std_ulogic; y: out std_ulogic);
    end component;

end apkg;
