package std is end;
