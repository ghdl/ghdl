entity t1 is
	err;
end t1;
