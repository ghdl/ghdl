entity ent is
end entity;

architecture a of ent is
    signal sig0 : integer_vector(0 to 7);
    signal sig1 : sig0'subtype(0 to 3);
begin
end;
