entity repro5 is
end;

architecture behav of repro5 is
  type states_t is (s0, s1, s2);
begin
end behav;
