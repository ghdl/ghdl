library ieee;use ieee.std_logic_1164;entity ghdlcrash is
port(a:std'u);end ghdlcrash;architecture h of g is--
function m(a:n)return l is
variable m:u;begin--
end function;begin
end architecture;