entity c is end entity;
architecture d of c is
signal foo: bit;
begin
foo <= '1';
end d;
