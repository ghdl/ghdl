package a is
end package a;
