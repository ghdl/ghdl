package cst is
  function four return natural;
end cst;

package body cst is
  function four return natural is
  begin
    return 4;
  end four;
end cst;
