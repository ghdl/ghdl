
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc224.vhd,v 1.2 2001-10-26 16:30:16 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c03s01b01x00p07n01i00224ent IS
END c03s01b01x00p07n01i00224ent;

ARCHITECTURE c03s01b01x00p07n01i00224arch OF c03s01b01x00p07n01i00224ent IS
  type ENUM1 is (FF, GG);
  type ENUM2 is (GG, HH);
  type ENUM3 is (FALSE);
  type ENUM4 is ('A', 'Z');
BEGIN
  TESTING: PROCESS
  BEGIN
    if ('A' = 'Z') then
      k := 5;
    end if;
    assert NOT( k=5 )
      report "***PASSED TEST: c03s01b01x00p07n01i00224"
      severity NOTE;
    assert ( k=5 )
      report "***FAILED TEST: c03s01b01x00p07n01i00224 - Literal cannot be determined." 
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c03s01b01x00p07n01i00224arch;
