entity compon is
end;

architecture behav of compon is
  signal s : bit;
begin
  inst: unknown
    port map (s => s);
end behav;
