�� - -   T h i s   i s   u t f - 1 6   B E   e n c o d i n g ,   w i t h   a   B O M . 
 
 p a c k a g e   p 1   i s 
 e n d   p 1 ; 
 
