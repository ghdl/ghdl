library ieee;
use ieee.std_logic_textio;

entity tb is
end tb;
