
-- Copyright (C) 2001 Bill Billowitch.

-- Some of the work to develop this test suite was done with Air Force
-- support.  The Air Force and Bill Billowitch assume no
-- responsibilities for this software.

-- This file is part of VESTs (Vhdl tESTs).

-- VESTs is free software; you can redistribute it and/or modify it
-- under the terms of the GNU General Public License as published by the
-- Free Software Foundation; either version 2 of the License, or (at
-- your option) any later version. 

-- VESTs is distributed in the hope that it will be useful, but WITHOUT
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
-- FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
-- for more details. 

-- You should have received a copy of the GNU General Public License
-- along with VESTs; if not, write to the Free Software Foundation,
-- Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 

-- ---------------------------------------------------------------------
--
-- $Id: tc2690.vhd,v 1.2 2001-10-26 16:29:49 paw Exp $
-- $Revision: 1.2 $
--
-- ---------------------------------------------------------------------

ENTITY c13s04b01x00p02n01i02690ent IS
  constant TIP_OFTHEICE    : Integer := 10 ;
  constant TIPOFTHEICE     : Real    := 0.546 ;
  constant T1       : Real := 3.14159_26 ;
  constant T2       : Real := 1.0E+6 ; --- No_failure_here
END c13s04b01x00p02n01i02690ent;

ARCHITECTURE c13s04b01x00p02n01i02690arch OF c13s04b01x00p02n01i02690ent IS

BEGIN
  TESTING: PROCESS
  BEGIN
    assert NOT(   TIP_OFTHEICE = 10   and
                  TIPOFTHEICE  = 0.546   and
                  T1        =3.14159_26   and
                  T2        = 1.0E+6   )
      report "***PASSED TEST: c13s04b01x00p02n01i02690"
      severity NOTE;
    assert (   TIP_OFTHEICE = 10   and
               TIPOFTHEICE  = 0.546   and
               T1        =3.14159_26   and
               T2        = 1.0E+6   )
      report "***FAILED TEST: c13s04b01x00p02n01i02690 - Correct decimal literal test failed."
      severity ERROR;
    wait;
  END PROCESS TESTING;

END c13s04b01x00p02n01i02690arch;
