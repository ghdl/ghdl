library ieee;
use ieee.std_logic_1164.all;

entity bug is
end bug;

architecture behavior of bug is
begin
    var1 : std_logic(1 downto 0);
end behavior;
