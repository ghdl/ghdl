package p is
  type rec is record
    a : bit; --  Comment for :a:
    b : bit; --  For :b:
  end record;
end p;
